module STI8_R5_23331543(in,out);
  input[15:0] in;
  output out;
  reg out;
  always@(in)
  begin
    case(in)
   0: out<=0;
   1: out<=0;
   2: out<=0;
   3: out<=0;
   4: out<=1;
   5: out<=0;
   6: out<=0;
   7: out<=1;
   8: out<=0;
   9: out<=1;
   10: out<=0;
   11: out<=1;
   12: out<=1;
   13: out<=1;
   14: out<=0;
   15: out<=0;
   16: out<=1;
   17: out<=1;
   18: out<=1;
   19: out<=1;
   20: out<=0;
   21: out<=1;
   22: out<=1;
   23: out<=0;
   24: out<=1;
   25: out<=0;
   26: out<=1;
   27: out<=0;
   28: out<=0;
   29: out<=0;
   30: out<=1;
   31: out<=1;
   32: out<=0;
   33: out<=0;
   34: out<=0;
   35: out<=0;
   36: out<=1;
   37: out<=0;
   38: out<=0;
   39: out<=1;
   40: out<=0;
   41: out<=1;
   42: out<=0;
   43: out<=1;
   44: out<=1;
   45: out<=1;
   46: out<=0;
   47: out<=0;
   48: out<=1;
   49: out<=1;
   50: out<=1;
   51: out<=1;
   52: out<=0;
   53: out<=1;
   54: out<=1;
   55: out<=0;
   56: out<=1;
   57: out<=0;
   58: out<=1;
   59: out<=0;
   60: out<=0;
   61: out<=0;
   62: out<=1;
   63: out<=1;
   64: out<=1;
   65: out<=1;
   66: out<=1;
   67: out<=1;
   68: out<=0;
   69: out<=1;
   70: out<=1;
   71: out<=0;
   72: out<=1;
   73: out<=0;
   74: out<=1;
   75: out<=0;
   76: out<=0;
   77: out<=0;
   78: out<=1;
   79: out<=1;
   80: out<=1;
   81: out<=1;
   82: out<=1;
   83: out<=1;
   84: out<=0;
   85: out<=1;
   86: out<=1;
   87: out<=0;
   88: out<=1;
   89: out<=0;
   90: out<=1;
   91: out<=0;
   92: out<=0;
   93: out<=0;
   94: out<=1;
   95: out<=1;
   96: out<=0;
   97: out<=0;
   98: out<=0;
   99: out<=0;
   100: out<=1;
   101: out<=0;
   102: out<=0;
   103: out<=1;
   104: out<=0;
   105: out<=1;
   106: out<=0;
   107: out<=1;
   108: out<=1;
   109: out<=1;
   110: out<=0;
   111: out<=0;
   112: out<=0;
   113: out<=0;
   114: out<=0;
   115: out<=0;
   116: out<=1;
   117: out<=0;
   118: out<=0;
   119: out<=1;
   120: out<=0;
   121: out<=1;
   122: out<=0;
   123: out<=1;
   124: out<=1;
   125: out<=1;
   126: out<=0;
   127: out<=0;
   128: out<=0;
   129: out<=0;
   130: out<=0;
   131: out<=0;
   132: out<=1;
   133: out<=0;
   134: out<=0;
   135: out<=1;
   136: out<=0;
   137: out<=1;
   138: out<=0;
   139: out<=1;
   140: out<=1;
   141: out<=1;
   142: out<=0;
   143: out<=0;
   144: out<=0;
   145: out<=0;
   146: out<=0;
   147: out<=0;
   148: out<=1;
   149: out<=0;
   150: out<=0;
   151: out<=1;
   152: out<=0;
   153: out<=1;
   154: out<=0;
   155: out<=1;
   156: out<=1;
   157: out<=1;
   158: out<=0;
   159: out<=0;
   160: out<=0;
   161: out<=0;
   162: out<=0;
   163: out<=0;
   164: out<=1;
   165: out<=0;
   166: out<=0;
   167: out<=1;
   168: out<=0;
   169: out<=1;
   170: out<=0;
   171: out<=1;
   172: out<=1;
   173: out<=1;
   174: out<=0;
   175: out<=0;
   176: out<=0;
   177: out<=0;
   178: out<=0;
   179: out<=0;
   180: out<=1;
   181: out<=0;
   182: out<=0;
   183: out<=1;
   184: out<=0;
   185: out<=1;
   186: out<=0;
   187: out<=1;
   188: out<=1;
   189: out<=1;
   190: out<=0;
   191: out<=0;
   192: out<=1;
   193: out<=1;
   194: out<=1;
   195: out<=1;
   196: out<=0;
   197: out<=1;
   198: out<=1;
   199: out<=0;
   200: out<=1;
   201: out<=0;
   202: out<=1;
   203: out<=0;
   204: out<=0;
   205: out<=0;
   206: out<=1;
   207: out<=1;
   208: out<=0;
   209: out<=0;
   210: out<=0;
   211: out<=0;
   212: out<=1;
   213: out<=0;
   214: out<=0;
   215: out<=1;
   216: out<=0;
   217: out<=1;
   218: out<=0;
   219: out<=1;
   220: out<=1;
   221: out<=1;
   222: out<=0;
   223: out<=0;
   224: out<=0;
   225: out<=0;
   226: out<=0;
   227: out<=0;
   228: out<=1;
   229: out<=0;
   230: out<=0;
   231: out<=1;
   232: out<=0;
   233: out<=1;
   234: out<=0;
   235: out<=1;
   236: out<=1;
   237: out<=1;
   238: out<=0;
   239: out<=0;
   240: out<=1;
   241: out<=1;
   242: out<=1;
   243: out<=1;
   244: out<=0;
   245: out<=1;
   246: out<=1;
   247: out<=0;
   248: out<=1;
   249: out<=0;
   250: out<=1;
   251: out<=0;
   252: out<=0;
   253: out<=0;
   254: out<=1;
   255: out<=1;
   256: out<=0;
   257: out<=1;
   258: out<=1;
   259: out<=0;
   260: out<=0;
   261: out<=0;
   262: out<=0;
   263: out<=0;
   264: out<=1;
   265: out<=1;
   266: out<=0;
   267: out<=0;
   268: out<=1;
   269: out<=0;
   270: out<=1;
   271: out<=0;
   272: out<=0;
   273: out<=1;
   274: out<=1;
   275: out<=0;
   276: out<=0;
   277: out<=0;
   278: out<=0;
   279: out<=0;
   280: out<=1;
   281: out<=1;
   282: out<=0;
   283: out<=0;
   284: out<=1;
   285: out<=0;
   286: out<=1;
   287: out<=0;
   288: out<=1;
   289: out<=0;
   290: out<=0;
   291: out<=1;
   292: out<=1;
   293: out<=1;
   294: out<=1;
   295: out<=1;
   296: out<=0;
   297: out<=0;
   298: out<=1;
   299: out<=1;
   300: out<=0;
   301: out<=1;
   302: out<=0;
   303: out<=1;
   304: out<=1;
   305: out<=0;
   306: out<=0;
   307: out<=1;
   308: out<=1;
   309: out<=1;
   310: out<=1;
   311: out<=1;
   312: out<=0;
   313: out<=0;
   314: out<=1;
   315: out<=1;
   316: out<=0;
   317: out<=1;
   318: out<=0;
   319: out<=1;
   320: out<=1;
   321: out<=0;
   322: out<=0;
   323: out<=1;
   324: out<=1;
   325: out<=1;
   326: out<=1;
   327: out<=1;
   328: out<=0;
   329: out<=0;
   330: out<=1;
   331: out<=1;
   332: out<=0;
   333: out<=1;
   334: out<=0;
   335: out<=1;
   336: out<=0;
   337: out<=1;
   338: out<=1;
   339: out<=0;
   340: out<=0;
   341: out<=0;
   342: out<=0;
   343: out<=0;
   344: out<=1;
   345: out<=1;
   346: out<=0;
   347: out<=0;
   348: out<=1;
   349: out<=0;
   350: out<=1;
   351: out<=0;
   352: out<=1;
   353: out<=0;
   354: out<=0;
   355: out<=1;
   356: out<=1;
   357: out<=1;
   358: out<=1;
   359: out<=1;
   360: out<=0;
   361: out<=0;
   362: out<=1;
   363: out<=1;
   364: out<=0;
   365: out<=1;
   366: out<=0;
   367: out<=1;
   368: out<=0;
   369: out<=1;
   370: out<=1;
   371: out<=0;
   372: out<=0;
   373: out<=0;
   374: out<=0;
   375: out<=0;
   376: out<=1;
   377: out<=1;
   378: out<=0;
   379: out<=0;
   380: out<=1;
   381: out<=0;
   382: out<=1;
   383: out<=0;
   384: out<=0;
   385: out<=1;
   386: out<=1;
   387: out<=0;
   388: out<=0;
   389: out<=0;
   390: out<=0;
   391: out<=0;
   392: out<=1;
   393: out<=1;
   394: out<=0;
   395: out<=0;
   396: out<=1;
   397: out<=0;
   398: out<=1;
   399: out<=0;
   400: out<=1;
   401: out<=0;
   402: out<=0;
   403: out<=1;
   404: out<=1;
   405: out<=1;
   406: out<=1;
   407: out<=1;
   408: out<=0;
   409: out<=0;
   410: out<=1;
   411: out<=1;
   412: out<=0;
   413: out<=1;
   414: out<=0;
   415: out<=1;
   416: out<=1;
   417: out<=0;
   418: out<=0;
   419: out<=1;
   420: out<=1;
   421: out<=1;
   422: out<=1;
   423: out<=1;
   424: out<=0;
   425: out<=0;
   426: out<=1;
   427: out<=1;
   428: out<=0;
   429: out<=1;
   430: out<=0;
   431: out<=1;
   432: out<=0;
   433: out<=1;
   434: out<=1;
   435: out<=0;
   436: out<=0;
   437: out<=0;
   438: out<=0;
   439: out<=0;
   440: out<=1;
   441: out<=1;
   442: out<=0;
   443: out<=0;
   444: out<=1;
   445: out<=0;
   446: out<=1;
   447: out<=0;
   448: out<=1;
   449: out<=0;
   450: out<=0;
   451: out<=1;
   452: out<=1;
   453: out<=1;
   454: out<=1;
   455: out<=1;
   456: out<=0;
   457: out<=0;
   458: out<=1;
   459: out<=1;
   460: out<=0;
   461: out<=1;
   462: out<=0;
   463: out<=1;
   464: out<=1;
   465: out<=0;
   466: out<=0;
   467: out<=1;
   468: out<=1;
   469: out<=1;
   470: out<=1;
   471: out<=1;
   472: out<=0;
   473: out<=0;
   474: out<=1;
   475: out<=1;
   476: out<=0;
   477: out<=1;
   478: out<=0;
   479: out<=1;
   480: out<=1;
   481: out<=0;
   482: out<=0;
   483: out<=1;
   484: out<=1;
   485: out<=1;
   486: out<=1;
   487: out<=1;
   488: out<=0;
   489: out<=0;
   490: out<=1;
   491: out<=1;
   492: out<=0;
   493: out<=1;
   494: out<=0;
   495: out<=1;
   496: out<=1;
   497: out<=0;
   498: out<=0;
   499: out<=1;
   500: out<=1;
   501: out<=1;
   502: out<=1;
   503: out<=1;
   504: out<=0;
   505: out<=0;
   506: out<=1;
   507: out<=1;
   508: out<=0;
   509: out<=1;
   510: out<=0;
   511: out<=1;
   512: out<=0;
   513: out<=1;
   514: out<=0;
   515: out<=1;
   516: out<=0;
   517: out<=0;
   518: out<=1;
   519: out<=1;
   520: out<=0;
   521: out<=0;
   522: out<=0;
   523: out<=0;
   524: out<=0;
   525: out<=1;
   526: out<=1;
   527: out<=0;
   528: out<=0;
   529: out<=1;
   530: out<=0;
   531: out<=1;
   532: out<=0;
   533: out<=0;
   534: out<=1;
   535: out<=1;
   536: out<=0;
   537: out<=0;
   538: out<=0;
   539: out<=0;
   540: out<=0;
   541: out<=1;
   542: out<=1;
   543: out<=0;
   544: out<=0;
   545: out<=1;
   546: out<=0;
   547: out<=1;
   548: out<=0;
   549: out<=0;
   550: out<=1;
   551: out<=1;
   552: out<=0;
   553: out<=0;
   554: out<=0;
   555: out<=0;
   556: out<=0;
   557: out<=1;
   558: out<=1;
   559: out<=0;
   560: out<=0;
   561: out<=1;
   562: out<=0;
   563: out<=1;
   564: out<=0;
   565: out<=0;
   566: out<=1;
   567: out<=1;
   568: out<=0;
   569: out<=0;
   570: out<=0;
   571: out<=0;
   572: out<=0;
   573: out<=1;
   574: out<=1;
   575: out<=0;
   576: out<=1;
   577: out<=0;
   578: out<=1;
   579: out<=0;
   580: out<=1;
   581: out<=1;
   582: out<=0;
   583: out<=0;
   584: out<=1;
   585: out<=1;
   586: out<=1;
   587: out<=1;
   588: out<=1;
   589: out<=0;
   590: out<=0;
   591: out<=1;
   592: out<=0;
   593: out<=1;
   594: out<=0;
   595: out<=1;
   596: out<=0;
   597: out<=0;
   598: out<=1;
   599: out<=1;
   600: out<=0;
   601: out<=0;
   602: out<=0;
   603: out<=0;
   604: out<=0;
   605: out<=1;
   606: out<=1;
   607: out<=0;
   608: out<=0;
   609: out<=1;
   610: out<=0;
   611: out<=1;
   612: out<=0;
   613: out<=0;
   614: out<=1;
   615: out<=1;
   616: out<=0;
   617: out<=0;
   618: out<=0;
   619: out<=0;
   620: out<=0;
   621: out<=1;
   622: out<=1;
   623: out<=0;
   624: out<=1;
   625: out<=0;
   626: out<=1;
   627: out<=0;
   628: out<=1;
   629: out<=1;
   630: out<=0;
   631: out<=0;
   632: out<=1;
   633: out<=1;
   634: out<=1;
   635: out<=1;
   636: out<=1;
   637: out<=0;
   638: out<=0;
   639: out<=1;
   640: out<=0;
   641: out<=1;
   642: out<=0;
   643: out<=1;
   644: out<=0;
   645: out<=0;
   646: out<=1;
   647: out<=1;
   648: out<=0;
   649: out<=0;
   650: out<=0;
   651: out<=0;
   652: out<=0;
   653: out<=1;
   654: out<=1;
   655: out<=0;
   656: out<=1;
   657: out<=0;
   658: out<=1;
   659: out<=0;
   660: out<=1;
   661: out<=1;
   662: out<=0;
   663: out<=0;
   664: out<=1;
   665: out<=1;
   666: out<=1;
   667: out<=1;
   668: out<=1;
   669: out<=0;
   670: out<=0;
   671: out<=1;
   672: out<=0;
   673: out<=1;
   674: out<=0;
   675: out<=1;
   676: out<=0;
   677: out<=0;
   678: out<=1;
   679: out<=1;
   680: out<=0;
   681: out<=0;
   682: out<=0;
   683: out<=0;
   684: out<=0;
   685: out<=1;
   686: out<=1;
   687: out<=0;
   688: out<=1;
   689: out<=0;
   690: out<=1;
   691: out<=0;
   692: out<=1;
   693: out<=1;
   694: out<=0;
   695: out<=0;
   696: out<=1;
   697: out<=1;
   698: out<=1;
   699: out<=1;
   700: out<=1;
   701: out<=0;
   702: out<=0;
   703: out<=1;
   704: out<=1;
   705: out<=0;
   706: out<=1;
   707: out<=0;
   708: out<=1;
   709: out<=1;
   710: out<=0;
   711: out<=0;
   712: out<=1;
   713: out<=1;
   714: out<=1;
   715: out<=1;
   716: out<=1;
   717: out<=0;
   718: out<=0;
   719: out<=1;
   720: out<=1;
   721: out<=0;
   722: out<=1;
   723: out<=0;
   724: out<=1;
   725: out<=1;
   726: out<=0;
   727: out<=0;
   728: out<=1;
   729: out<=1;
   730: out<=1;
   731: out<=1;
   732: out<=1;
   733: out<=0;
   734: out<=0;
   735: out<=1;
   736: out<=0;
   737: out<=1;
   738: out<=0;
   739: out<=1;
   740: out<=0;
   741: out<=0;
   742: out<=1;
   743: out<=1;
   744: out<=0;
   745: out<=0;
   746: out<=0;
   747: out<=0;
   748: out<=0;
   749: out<=1;
   750: out<=1;
   751: out<=0;
   752: out<=0;
   753: out<=1;
   754: out<=0;
   755: out<=1;
   756: out<=0;
   757: out<=0;
   758: out<=1;
   759: out<=1;
   760: out<=0;
   761: out<=0;
   762: out<=0;
   763: out<=0;
   764: out<=0;
   765: out<=1;
   766: out<=1;
   767: out<=0;
   768: out<=0;
   769: out<=0;
   770: out<=1;
   771: out<=1;
   772: out<=1;
   773: out<=0;
   774: out<=1;
   775: out<=0;
   776: out<=1;
   777: out<=0;
   778: out<=0;
   779: out<=1;
   780: out<=0;
   781: out<=0;
   782: out<=0;
   783: out<=0;
   784: out<=1;
   785: out<=1;
   786: out<=0;
   787: out<=0;
   788: out<=0;
   789: out<=1;
   790: out<=0;
   791: out<=1;
   792: out<=0;
   793: out<=1;
   794: out<=1;
   795: out<=0;
   796: out<=1;
   797: out<=1;
   798: out<=1;
   799: out<=1;
   800: out<=1;
   801: out<=1;
   802: out<=0;
   803: out<=0;
   804: out<=0;
   805: out<=1;
   806: out<=0;
   807: out<=1;
   808: out<=0;
   809: out<=1;
   810: out<=1;
   811: out<=0;
   812: out<=1;
   813: out<=1;
   814: out<=1;
   815: out<=1;
   816: out<=0;
   817: out<=0;
   818: out<=1;
   819: out<=1;
   820: out<=1;
   821: out<=0;
   822: out<=1;
   823: out<=0;
   824: out<=1;
   825: out<=0;
   826: out<=0;
   827: out<=1;
   828: out<=0;
   829: out<=0;
   830: out<=0;
   831: out<=0;
   832: out<=1;
   833: out<=1;
   834: out<=0;
   835: out<=0;
   836: out<=0;
   837: out<=1;
   838: out<=0;
   839: out<=1;
   840: out<=0;
   841: out<=1;
   842: out<=1;
   843: out<=0;
   844: out<=1;
   845: out<=1;
   846: out<=1;
   847: out<=1;
   848: out<=1;
   849: out<=1;
   850: out<=0;
   851: out<=0;
   852: out<=0;
   853: out<=1;
   854: out<=0;
   855: out<=1;
   856: out<=0;
   857: out<=1;
   858: out<=1;
   859: out<=0;
   860: out<=1;
   861: out<=1;
   862: out<=1;
   863: out<=1;
   864: out<=1;
   865: out<=1;
   866: out<=0;
   867: out<=0;
   868: out<=0;
   869: out<=1;
   870: out<=0;
   871: out<=1;
   872: out<=0;
   873: out<=1;
   874: out<=1;
   875: out<=0;
   876: out<=1;
   877: out<=1;
   878: out<=1;
   879: out<=1;
   880: out<=1;
   881: out<=1;
   882: out<=0;
   883: out<=0;
   884: out<=0;
   885: out<=1;
   886: out<=0;
   887: out<=1;
   888: out<=0;
   889: out<=1;
   890: out<=1;
   891: out<=0;
   892: out<=1;
   893: out<=1;
   894: out<=1;
   895: out<=1;
   896: out<=0;
   897: out<=0;
   898: out<=1;
   899: out<=1;
   900: out<=1;
   901: out<=0;
   902: out<=1;
   903: out<=0;
   904: out<=1;
   905: out<=0;
   906: out<=0;
   907: out<=1;
   908: out<=0;
   909: out<=0;
   910: out<=0;
   911: out<=0;
   912: out<=0;
   913: out<=0;
   914: out<=1;
   915: out<=1;
   916: out<=1;
   917: out<=0;
   918: out<=1;
   919: out<=0;
   920: out<=1;
   921: out<=0;
   922: out<=0;
   923: out<=1;
   924: out<=0;
   925: out<=0;
   926: out<=0;
   927: out<=0;
   928: out<=1;
   929: out<=1;
   930: out<=0;
   931: out<=0;
   932: out<=0;
   933: out<=1;
   934: out<=0;
   935: out<=1;
   936: out<=0;
   937: out<=1;
   938: out<=1;
   939: out<=0;
   940: out<=1;
   941: out<=1;
   942: out<=1;
   943: out<=1;
   944: out<=1;
   945: out<=1;
   946: out<=0;
   947: out<=0;
   948: out<=0;
   949: out<=1;
   950: out<=0;
   951: out<=1;
   952: out<=0;
   953: out<=1;
   954: out<=1;
   955: out<=0;
   956: out<=1;
   957: out<=1;
   958: out<=1;
   959: out<=1;
   960: out<=1;
   961: out<=1;
   962: out<=0;
   963: out<=0;
   964: out<=0;
   965: out<=1;
   966: out<=0;
   967: out<=1;
   968: out<=0;
   969: out<=1;
   970: out<=1;
   971: out<=0;
   972: out<=1;
   973: out<=1;
   974: out<=1;
   975: out<=1;
   976: out<=0;
   977: out<=0;
   978: out<=1;
   979: out<=1;
   980: out<=1;
   981: out<=0;
   982: out<=1;
   983: out<=0;
   984: out<=1;
   985: out<=0;
   986: out<=0;
   987: out<=1;
   988: out<=0;
   989: out<=0;
   990: out<=0;
   991: out<=0;
   992: out<=1;
   993: out<=1;
   994: out<=0;
   995: out<=0;
   996: out<=0;
   997: out<=1;
   998: out<=0;
   999: out<=1;
   1000: out<=0;
   1001: out<=1;
   1002: out<=1;
   1003: out<=0;
   1004: out<=1;
   1005: out<=1;
   1006: out<=1;
   1007: out<=1;
   1008: out<=0;
   1009: out<=0;
   1010: out<=1;
   1011: out<=1;
   1012: out<=1;
   1013: out<=0;
   1014: out<=1;
   1015: out<=0;
   1016: out<=1;
   1017: out<=0;
   1018: out<=0;
   1019: out<=1;
   1020: out<=0;
   1021: out<=0;
   1022: out<=0;
   1023: out<=0;
   1024: out<=0;
   1025: out<=1;
   1026: out<=1;
   1027: out<=0;
   1028: out<=1;
   1029: out<=1;
   1030: out<=1;
   1031: out<=1;
   1032: out<=0;
   1033: out<=0;
   1034: out<=1;
   1035: out<=1;
   1036: out<=1;
   1037: out<=0;
   1038: out<=1;
   1039: out<=0;
   1040: out<=1;
   1041: out<=0;
   1042: out<=0;
   1043: out<=1;
   1044: out<=0;
   1045: out<=0;
   1046: out<=0;
   1047: out<=0;
   1048: out<=1;
   1049: out<=1;
   1050: out<=0;
   1051: out<=0;
   1052: out<=0;
   1053: out<=1;
   1054: out<=0;
   1055: out<=1;
   1056: out<=0;
   1057: out<=1;
   1058: out<=1;
   1059: out<=0;
   1060: out<=1;
   1061: out<=1;
   1062: out<=1;
   1063: out<=1;
   1064: out<=0;
   1065: out<=0;
   1066: out<=1;
   1067: out<=1;
   1068: out<=1;
   1069: out<=0;
   1070: out<=1;
   1071: out<=0;
   1072: out<=1;
   1073: out<=0;
   1074: out<=0;
   1075: out<=1;
   1076: out<=0;
   1077: out<=0;
   1078: out<=0;
   1079: out<=0;
   1080: out<=1;
   1081: out<=1;
   1082: out<=0;
   1083: out<=0;
   1084: out<=0;
   1085: out<=1;
   1086: out<=0;
   1087: out<=1;
   1088: out<=1;
   1089: out<=0;
   1090: out<=0;
   1091: out<=1;
   1092: out<=0;
   1093: out<=0;
   1094: out<=0;
   1095: out<=0;
   1096: out<=1;
   1097: out<=1;
   1098: out<=0;
   1099: out<=0;
   1100: out<=0;
   1101: out<=1;
   1102: out<=0;
   1103: out<=1;
   1104: out<=1;
   1105: out<=0;
   1106: out<=0;
   1107: out<=1;
   1108: out<=0;
   1109: out<=0;
   1110: out<=0;
   1111: out<=0;
   1112: out<=1;
   1113: out<=1;
   1114: out<=0;
   1115: out<=0;
   1116: out<=0;
   1117: out<=1;
   1118: out<=0;
   1119: out<=1;
   1120: out<=0;
   1121: out<=1;
   1122: out<=1;
   1123: out<=0;
   1124: out<=1;
   1125: out<=1;
   1126: out<=1;
   1127: out<=1;
   1128: out<=0;
   1129: out<=0;
   1130: out<=1;
   1131: out<=1;
   1132: out<=1;
   1133: out<=0;
   1134: out<=1;
   1135: out<=0;
   1136: out<=0;
   1137: out<=1;
   1138: out<=1;
   1139: out<=0;
   1140: out<=1;
   1141: out<=1;
   1142: out<=1;
   1143: out<=1;
   1144: out<=0;
   1145: out<=0;
   1146: out<=1;
   1147: out<=1;
   1148: out<=1;
   1149: out<=0;
   1150: out<=1;
   1151: out<=0;
   1152: out<=0;
   1153: out<=1;
   1154: out<=1;
   1155: out<=0;
   1156: out<=1;
   1157: out<=1;
   1158: out<=1;
   1159: out<=1;
   1160: out<=0;
   1161: out<=0;
   1162: out<=1;
   1163: out<=1;
   1164: out<=1;
   1165: out<=0;
   1166: out<=1;
   1167: out<=0;
   1168: out<=0;
   1169: out<=1;
   1170: out<=1;
   1171: out<=0;
   1172: out<=1;
   1173: out<=1;
   1174: out<=1;
   1175: out<=1;
   1176: out<=0;
   1177: out<=0;
   1178: out<=1;
   1179: out<=1;
   1180: out<=1;
   1181: out<=0;
   1182: out<=1;
   1183: out<=0;
   1184: out<=0;
   1185: out<=1;
   1186: out<=1;
   1187: out<=0;
   1188: out<=1;
   1189: out<=1;
   1190: out<=1;
   1191: out<=1;
   1192: out<=0;
   1193: out<=0;
   1194: out<=1;
   1195: out<=1;
   1196: out<=1;
   1197: out<=0;
   1198: out<=1;
   1199: out<=0;
   1200: out<=0;
   1201: out<=1;
   1202: out<=1;
   1203: out<=0;
   1204: out<=1;
   1205: out<=1;
   1206: out<=1;
   1207: out<=1;
   1208: out<=0;
   1209: out<=0;
   1210: out<=1;
   1211: out<=1;
   1212: out<=1;
   1213: out<=0;
   1214: out<=1;
   1215: out<=0;
   1216: out<=1;
   1217: out<=0;
   1218: out<=0;
   1219: out<=1;
   1220: out<=0;
   1221: out<=0;
   1222: out<=0;
   1223: out<=0;
   1224: out<=1;
   1225: out<=1;
   1226: out<=0;
   1227: out<=0;
   1228: out<=0;
   1229: out<=1;
   1230: out<=0;
   1231: out<=1;
   1232: out<=0;
   1233: out<=1;
   1234: out<=1;
   1235: out<=0;
   1236: out<=1;
   1237: out<=1;
   1238: out<=1;
   1239: out<=1;
   1240: out<=0;
   1241: out<=0;
   1242: out<=1;
   1243: out<=1;
   1244: out<=1;
   1245: out<=0;
   1246: out<=1;
   1247: out<=0;
   1248: out<=0;
   1249: out<=1;
   1250: out<=1;
   1251: out<=0;
   1252: out<=1;
   1253: out<=1;
   1254: out<=1;
   1255: out<=1;
   1256: out<=0;
   1257: out<=0;
   1258: out<=1;
   1259: out<=1;
   1260: out<=1;
   1261: out<=0;
   1262: out<=1;
   1263: out<=0;
   1264: out<=1;
   1265: out<=0;
   1266: out<=0;
   1267: out<=1;
   1268: out<=0;
   1269: out<=0;
   1270: out<=0;
   1271: out<=0;
   1272: out<=1;
   1273: out<=1;
   1274: out<=0;
   1275: out<=0;
   1276: out<=0;
   1277: out<=1;
   1278: out<=0;
   1279: out<=1;
   1280: out<=1;
   1281: out<=1;
   1282: out<=1;
   1283: out<=1;
   1284: out<=1;
   1285: out<=0;
   1286: out<=0;
   1287: out<=1;
   1288: out<=0;
   1289: out<=1;
   1290: out<=0;
   1291: out<=1;
   1292: out<=0;
   1293: out<=0;
   1294: out<=1;
   1295: out<=1;
   1296: out<=1;
   1297: out<=1;
   1298: out<=1;
   1299: out<=1;
   1300: out<=1;
   1301: out<=0;
   1302: out<=0;
   1303: out<=1;
   1304: out<=0;
   1305: out<=1;
   1306: out<=0;
   1307: out<=1;
   1308: out<=0;
   1309: out<=0;
   1310: out<=1;
   1311: out<=1;
   1312: out<=0;
   1313: out<=0;
   1314: out<=0;
   1315: out<=0;
   1316: out<=0;
   1317: out<=1;
   1318: out<=1;
   1319: out<=0;
   1320: out<=1;
   1321: out<=0;
   1322: out<=1;
   1323: out<=0;
   1324: out<=1;
   1325: out<=1;
   1326: out<=0;
   1327: out<=0;
   1328: out<=0;
   1329: out<=0;
   1330: out<=0;
   1331: out<=0;
   1332: out<=0;
   1333: out<=1;
   1334: out<=1;
   1335: out<=0;
   1336: out<=1;
   1337: out<=0;
   1338: out<=1;
   1339: out<=0;
   1340: out<=1;
   1341: out<=1;
   1342: out<=0;
   1343: out<=0;
   1344: out<=0;
   1345: out<=0;
   1346: out<=0;
   1347: out<=0;
   1348: out<=0;
   1349: out<=1;
   1350: out<=1;
   1351: out<=0;
   1352: out<=1;
   1353: out<=0;
   1354: out<=1;
   1355: out<=0;
   1356: out<=1;
   1357: out<=1;
   1358: out<=0;
   1359: out<=0;
   1360: out<=1;
   1361: out<=1;
   1362: out<=1;
   1363: out<=1;
   1364: out<=1;
   1365: out<=0;
   1366: out<=0;
   1367: out<=1;
   1368: out<=0;
   1369: out<=1;
   1370: out<=0;
   1371: out<=1;
   1372: out<=0;
   1373: out<=0;
   1374: out<=1;
   1375: out<=1;
   1376: out<=0;
   1377: out<=0;
   1378: out<=0;
   1379: out<=0;
   1380: out<=0;
   1381: out<=1;
   1382: out<=1;
   1383: out<=0;
   1384: out<=1;
   1385: out<=0;
   1386: out<=1;
   1387: out<=0;
   1388: out<=1;
   1389: out<=1;
   1390: out<=0;
   1391: out<=0;
   1392: out<=1;
   1393: out<=1;
   1394: out<=1;
   1395: out<=1;
   1396: out<=1;
   1397: out<=0;
   1398: out<=0;
   1399: out<=1;
   1400: out<=0;
   1401: out<=1;
   1402: out<=0;
   1403: out<=1;
   1404: out<=0;
   1405: out<=0;
   1406: out<=1;
   1407: out<=1;
   1408: out<=1;
   1409: out<=1;
   1410: out<=1;
   1411: out<=1;
   1412: out<=1;
   1413: out<=0;
   1414: out<=0;
   1415: out<=1;
   1416: out<=0;
   1417: out<=1;
   1418: out<=0;
   1419: out<=1;
   1420: out<=0;
   1421: out<=0;
   1422: out<=1;
   1423: out<=1;
   1424: out<=0;
   1425: out<=0;
   1426: out<=0;
   1427: out<=0;
   1428: out<=0;
   1429: out<=1;
   1430: out<=1;
   1431: out<=0;
   1432: out<=1;
   1433: out<=0;
   1434: out<=1;
   1435: out<=0;
   1436: out<=1;
   1437: out<=1;
   1438: out<=0;
   1439: out<=0;
   1440: out<=0;
   1441: out<=0;
   1442: out<=0;
   1443: out<=0;
   1444: out<=0;
   1445: out<=1;
   1446: out<=1;
   1447: out<=0;
   1448: out<=1;
   1449: out<=0;
   1450: out<=1;
   1451: out<=0;
   1452: out<=1;
   1453: out<=1;
   1454: out<=0;
   1455: out<=0;
   1456: out<=1;
   1457: out<=1;
   1458: out<=1;
   1459: out<=1;
   1460: out<=1;
   1461: out<=0;
   1462: out<=0;
   1463: out<=1;
   1464: out<=0;
   1465: out<=1;
   1466: out<=0;
   1467: out<=1;
   1468: out<=0;
   1469: out<=0;
   1470: out<=1;
   1471: out<=1;
   1472: out<=0;
   1473: out<=0;
   1474: out<=0;
   1475: out<=0;
   1476: out<=0;
   1477: out<=1;
   1478: out<=1;
   1479: out<=0;
   1480: out<=1;
   1481: out<=0;
   1482: out<=1;
   1483: out<=0;
   1484: out<=1;
   1485: out<=1;
   1486: out<=0;
   1487: out<=0;
   1488: out<=0;
   1489: out<=0;
   1490: out<=0;
   1491: out<=0;
   1492: out<=0;
   1493: out<=1;
   1494: out<=1;
   1495: out<=0;
   1496: out<=1;
   1497: out<=0;
   1498: out<=1;
   1499: out<=0;
   1500: out<=1;
   1501: out<=1;
   1502: out<=0;
   1503: out<=0;
   1504: out<=0;
   1505: out<=0;
   1506: out<=0;
   1507: out<=0;
   1508: out<=0;
   1509: out<=1;
   1510: out<=1;
   1511: out<=0;
   1512: out<=1;
   1513: out<=0;
   1514: out<=1;
   1515: out<=0;
   1516: out<=1;
   1517: out<=1;
   1518: out<=0;
   1519: out<=0;
   1520: out<=0;
   1521: out<=0;
   1522: out<=0;
   1523: out<=0;
   1524: out<=0;
   1525: out<=1;
   1526: out<=1;
   1527: out<=0;
   1528: out<=1;
   1529: out<=0;
   1530: out<=1;
   1531: out<=0;
   1532: out<=1;
   1533: out<=1;
   1534: out<=0;
   1535: out<=0;
   1536: out<=1;
   1537: out<=1;
   1538: out<=0;
   1539: out<=0;
   1540: out<=1;
   1541: out<=0;
   1542: out<=1;
   1543: out<=0;
   1544: out<=1;
   1545: out<=0;
   1546: out<=0;
   1547: out<=1;
   1548: out<=1;
   1549: out<=1;
   1550: out<=1;
   1551: out<=1;
   1552: out<=1;
   1553: out<=1;
   1554: out<=0;
   1555: out<=0;
   1556: out<=1;
   1557: out<=0;
   1558: out<=1;
   1559: out<=0;
   1560: out<=1;
   1561: out<=0;
   1562: out<=0;
   1563: out<=1;
   1564: out<=1;
   1565: out<=1;
   1566: out<=1;
   1567: out<=1;
   1568: out<=1;
   1569: out<=1;
   1570: out<=0;
   1571: out<=0;
   1572: out<=1;
   1573: out<=0;
   1574: out<=1;
   1575: out<=0;
   1576: out<=1;
   1577: out<=0;
   1578: out<=0;
   1579: out<=1;
   1580: out<=1;
   1581: out<=1;
   1582: out<=1;
   1583: out<=1;
   1584: out<=1;
   1585: out<=1;
   1586: out<=0;
   1587: out<=0;
   1588: out<=1;
   1589: out<=0;
   1590: out<=1;
   1591: out<=0;
   1592: out<=1;
   1593: out<=0;
   1594: out<=0;
   1595: out<=1;
   1596: out<=1;
   1597: out<=1;
   1598: out<=1;
   1599: out<=1;
   1600: out<=0;
   1601: out<=0;
   1602: out<=1;
   1603: out<=1;
   1604: out<=0;
   1605: out<=1;
   1606: out<=0;
   1607: out<=1;
   1608: out<=0;
   1609: out<=1;
   1610: out<=1;
   1611: out<=0;
   1612: out<=0;
   1613: out<=0;
   1614: out<=0;
   1615: out<=0;
   1616: out<=1;
   1617: out<=1;
   1618: out<=0;
   1619: out<=0;
   1620: out<=1;
   1621: out<=0;
   1622: out<=1;
   1623: out<=0;
   1624: out<=1;
   1625: out<=0;
   1626: out<=0;
   1627: out<=1;
   1628: out<=1;
   1629: out<=1;
   1630: out<=1;
   1631: out<=1;
   1632: out<=1;
   1633: out<=1;
   1634: out<=0;
   1635: out<=0;
   1636: out<=1;
   1637: out<=0;
   1638: out<=1;
   1639: out<=0;
   1640: out<=1;
   1641: out<=0;
   1642: out<=0;
   1643: out<=1;
   1644: out<=1;
   1645: out<=1;
   1646: out<=1;
   1647: out<=1;
   1648: out<=0;
   1649: out<=0;
   1650: out<=1;
   1651: out<=1;
   1652: out<=0;
   1653: out<=1;
   1654: out<=0;
   1655: out<=1;
   1656: out<=0;
   1657: out<=1;
   1658: out<=1;
   1659: out<=0;
   1660: out<=0;
   1661: out<=0;
   1662: out<=0;
   1663: out<=0;
   1664: out<=1;
   1665: out<=1;
   1666: out<=0;
   1667: out<=0;
   1668: out<=1;
   1669: out<=0;
   1670: out<=1;
   1671: out<=0;
   1672: out<=1;
   1673: out<=0;
   1674: out<=0;
   1675: out<=1;
   1676: out<=1;
   1677: out<=1;
   1678: out<=1;
   1679: out<=1;
   1680: out<=0;
   1681: out<=0;
   1682: out<=1;
   1683: out<=1;
   1684: out<=0;
   1685: out<=1;
   1686: out<=0;
   1687: out<=1;
   1688: out<=0;
   1689: out<=1;
   1690: out<=1;
   1691: out<=0;
   1692: out<=0;
   1693: out<=0;
   1694: out<=0;
   1695: out<=0;
   1696: out<=1;
   1697: out<=1;
   1698: out<=0;
   1699: out<=0;
   1700: out<=1;
   1701: out<=0;
   1702: out<=1;
   1703: out<=0;
   1704: out<=1;
   1705: out<=0;
   1706: out<=0;
   1707: out<=1;
   1708: out<=1;
   1709: out<=1;
   1710: out<=1;
   1711: out<=1;
   1712: out<=0;
   1713: out<=0;
   1714: out<=1;
   1715: out<=1;
   1716: out<=0;
   1717: out<=1;
   1718: out<=0;
   1719: out<=1;
   1720: out<=0;
   1721: out<=1;
   1722: out<=1;
   1723: out<=0;
   1724: out<=0;
   1725: out<=0;
   1726: out<=0;
   1727: out<=0;
   1728: out<=0;
   1729: out<=0;
   1730: out<=1;
   1731: out<=1;
   1732: out<=0;
   1733: out<=1;
   1734: out<=0;
   1735: out<=1;
   1736: out<=0;
   1737: out<=1;
   1738: out<=1;
   1739: out<=0;
   1740: out<=0;
   1741: out<=0;
   1742: out<=0;
   1743: out<=0;
   1744: out<=0;
   1745: out<=0;
   1746: out<=1;
   1747: out<=1;
   1748: out<=0;
   1749: out<=1;
   1750: out<=0;
   1751: out<=1;
   1752: out<=0;
   1753: out<=1;
   1754: out<=1;
   1755: out<=0;
   1756: out<=0;
   1757: out<=0;
   1758: out<=0;
   1759: out<=0;
   1760: out<=1;
   1761: out<=1;
   1762: out<=0;
   1763: out<=0;
   1764: out<=1;
   1765: out<=0;
   1766: out<=1;
   1767: out<=0;
   1768: out<=1;
   1769: out<=0;
   1770: out<=0;
   1771: out<=1;
   1772: out<=1;
   1773: out<=1;
   1774: out<=1;
   1775: out<=1;
   1776: out<=1;
   1777: out<=1;
   1778: out<=0;
   1779: out<=0;
   1780: out<=1;
   1781: out<=0;
   1782: out<=1;
   1783: out<=0;
   1784: out<=1;
   1785: out<=0;
   1786: out<=0;
   1787: out<=1;
   1788: out<=1;
   1789: out<=1;
   1790: out<=1;
   1791: out<=1;
   1792: out<=0;
   1793: out<=1;
   1794: out<=0;
   1795: out<=1;
   1796: out<=1;
   1797: out<=1;
   1798: out<=0;
   1799: out<=0;
   1800: out<=1;
   1801: out<=1;
   1802: out<=1;
   1803: out<=1;
   1804: out<=0;
   1805: out<=1;
   1806: out<=1;
   1807: out<=0;
   1808: out<=1;
   1809: out<=0;
   1810: out<=1;
   1811: out<=0;
   1812: out<=0;
   1813: out<=0;
   1814: out<=1;
   1815: out<=1;
   1816: out<=0;
   1817: out<=0;
   1818: out<=0;
   1819: out<=0;
   1820: out<=1;
   1821: out<=0;
   1822: out<=0;
   1823: out<=1;
   1824: out<=1;
   1825: out<=0;
   1826: out<=1;
   1827: out<=0;
   1828: out<=0;
   1829: out<=0;
   1830: out<=1;
   1831: out<=1;
   1832: out<=0;
   1833: out<=0;
   1834: out<=0;
   1835: out<=0;
   1836: out<=1;
   1837: out<=0;
   1838: out<=0;
   1839: out<=1;
   1840: out<=0;
   1841: out<=1;
   1842: out<=0;
   1843: out<=1;
   1844: out<=1;
   1845: out<=1;
   1846: out<=0;
   1847: out<=0;
   1848: out<=1;
   1849: out<=1;
   1850: out<=1;
   1851: out<=1;
   1852: out<=0;
   1853: out<=1;
   1854: out<=1;
   1855: out<=0;
   1856: out<=1;
   1857: out<=0;
   1858: out<=1;
   1859: out<=0;
   1860: out<=0;
   1861: out<=0;
   1862: out<=1;
   1863: out<=1;
   1864: out<=0;
   1865: out<=0;
   1866: out<=0;
   1867: out<=0;
   1868: out<=1;
   1869: out<=0;
   1870: out<=0;
   1871: out<=1;
   1872: out<=1;
   1873: out<=0;
   1874: out<=1;
   1875: out<=0;
   1876: out<=0;
   1877: out<=0;
   1878: out<=1;
   1879: out<=1;
   1880: out<=0;
   1881: out<=0;
   1882: out<=0;
   1883: out<=0;
   1884: out<=1;
   1885: out<=0;
   1886: out<=0;
   1887: out<=1;
   1888: out<=1;
   1889: out<=0;
   1890: out<=1;
   1891: out<=0;
   1892: out<=0;
   1893: out<=0;
   1894: out<=1;
   1895: out<=1;
   1896: out<=0;
   1897: out<=0;
   1898: out<=0;
   1899: out<=0;
   1900: out<=1;
   1901: out<=0;
   1902: out<=0;
   1903: out<=1;
   1904: out<=1;
   1905: out<=0;
   1906: out<=1;
   1907: out<=0;
   1908: out<=0;
   1909: out<=0;
   1910: out<=1;
   1911: out<=1;
   1912: out<=0;
   1913: out<=0;
   1914: out<=0;
   1915: out<=0;
   1916: out<=1;
   1917: out<=0;
   1918: out<=0;
   1919: out<=1;
   1920: out<=0;
   1921: out<=1;
   1922: out<=0;
   1923: out<=1;
   1924: out<=1;
   1925: out<=1;
   1926: out<=0;
   1927: out<=0;
   1928: out<=1;
   1929: out<=1;
   1930: out<=1;
   1931: out<=1;
   1932: out<=0;
   1933: out<=1;
   1934: out<=1;
   1935: out<=0;
   1936: out<=0;
   1937: out<=1;
   1938: out<=0;
   1939: out<=1;
   1940: out<=1;
   1941: out<=1;
   1942: out<=0;
   1943: out<=0;
   1944: out<=1;
   1945: out<=1;
   1946: out<=1;
   1947: out<=1;
   1948: out<=0;
   1949: out<=1;
   1950: out<=1;
   1951: out<=0;
   1952: out<=1;
   1953: out<=0;
   1954: out<=1;
   1955: out<=0;
   1956: out<=0;
   1957: out<=0;
   1958: out<=1;
   1959: out<=1;
   1960: out<=0;
   1961: out<=0;
   1962: out<=0;
   1963: out<=0;
   1964: out<=1;
   1965: out<=0;
   1966: out<=0;
   1967: out<=1;
   1968: out<=1;
   1969: out<=0;
   1970: out<=1;
   1971: out<=0;
   1972: out<=0;
   1973: out<=0;
   1974: out<=1;
   1975: out<=1;
   1976: out<=0;
   1977: out<=0;
   1978: out<=0;
   1979: out<=0;
   1980: out<=1;
   1981: out<=0;
   1982: out<=0;
   1983: out<=1;
   1984: out<=1;
   1985: out<=0;
   1986: out<=1;
   1987: out<=0;
   1988: out<=0;
   1989: out<=0;
   1990: out<=1;
   1991: out<=1;
   1992: out<=0;
   1993: out<=0;
   1994: out<=0;
   1995: out<=0;
   1996: out<=1;
   1997: out<=0;
   1998: out<=0;
   1999: out<=1;
   2000: out<=0;
   2001: out<=1;
   2002: out<=0;
   2003: out<=1;
   2004: out<=1;
   2005: out<=1;
   2006: out<=0;
   2007: out<=0;
   2008: out<=1;
   2009: out<=1;
   2010: out<=1;
   2011: out<=1;
   2012: out<=0;
   2013: out<=1;
   2014: out<=1;
   2015: out<=0;
   2016: out<=1;
   2017: out<=0;
   2018: out<=1;
   2019: out<=0;
   2020: out<=0;
   2021: out<=0;
   2022: out<=1;
   2023: out<=1;
   2024: out<=0;
   2025: out<=0;
   2026: out<=0;
   2027: out<=0;
   2028: out<=1;
   2029: out<=0;
   2030: out<=0;
   2031: out<=1;
   2032: out<=0;
   2033: out<=1;
   2034: out<=0;
   2035: out<=1;
   2036: out<=1;
   2037: out<=1;
   2038: out<=0;
   2039: out<=0;
   2040: out<=1;
   2041: out<=1;
   2042: out<=1;
   2043: out<=1;
   2044: out<=0;
   2045: out<=1;
   2046: out<=1;
   2047: out<=0;
   2048: out<=0;
   2049: out<=1;
   2050: out<=0;
   2051: out<=1;
   2052: out<=1;
   2053: out<=1;
   2054: out<=0;
   2055: out<=0;
   2056: out<=0;
   2057: out<=0;
   2058: out<=0;
   2059: out<=0;
   2060: out<=1;
   2061: out<=0;
   2062: out<=0;
   2063: out<=1;
   2064: out<=1;
   2065: out<=0;
   2066: out<=1;
   2067: out<=0;
   2068: out<=0;
   2069: out<=0;
   2070: out<=1;
   2071: out<=1;
   2072: out<=1;
   2073: out<=1;
   2074: out<=1;
   2075: out<=1;
   2076: out<=0;
   2077: out<=1;
   2078: out<=1;
   2079: out<=0;
   2080: out<=0;
   2081: out<=1;
   2082: out<=0;
   2083: out<=1;
   2084: out<=1;
   2085: out<=1;
   2086: out<=0;
   2087: out<=0;
   2088: out<=0;
   2089: out<=0;
   2090: out<=0;
   2091: out<=0;
   2092: out<=1;
   2093: out<=0;
   2094: out<=0;
   2095: out<=1;
   2096: out<=1;
   2097: out<=0;
   2098: out<=1;
   2099: out<=0;
   2100: out<=0;
   2101: out<=0;
   2102: out<=1;
   2103: out<=1;
   2104: out<=1;
   2105: out<=1;
   2106: out<=1;
   2107: out<=1;
   2108: out<=0;
   2109: out<=1;
   2110: out<=1;
   2111: out<=0;
   2112: out<=1;
   2113: out<=0;
   2114: out<=1;
   2115: out<=0;
   2116: out<=0;
   2117: out<=0;
   2118: out<=1;
   2119: out<=1;
   2120: out<=1;
   2121: out<=1;
   2122: out<=1;
   2123: out<=1;
   2124: out<=0;
   2125: out<=1;
   2126: out<=1;
   2127: out<=0;
   2128: out<=1;
   2129: out<=0;
   2130: out<=1;
   2131: out<=0;
   2132: out<=0;
   2133: out<=0;
   2134: out<=1;
   2135: out<=1;
   2136: out<=1;
   2137: out<=1;
   2138: out<=1;
   2139: out<=1;
   2140: out<=0;
   2141: out<=1;
   2142: out<=1;
   2143: out<=0;
   2144: out<=0;
   2145: out<=1;
   2146: out<=0;
   2147: out<=1;
   2148: out<=1;
   2149: out<=1;
   2150: out<=0;
   2151: out<=0;
   2152: out<=0;
   2153: out<=0;
   2154: out<=0;
   2155: out<=0;
   2156: out<=1;
   2157: out<=0;
   2158: out<=0;
   2159: out<=1;
   2160: out<=0;
   2161: out<=1;
   2162: out<=0;
   2163: out<=1;
   2164: out<=1;
   2165: out<=1;
   2166: out<=0;
   2167: out<=0;
   2168: out<=0;
   2169: out<=0;
   2170: out<=0;
   2171: out<=0;
   2172: out<=1;
   2173: out<=0;
   2174: out<=0;
   2175: out<=1;
   2176: out<=0;
   2177: out<=1;
   2178: out<=0;
   2179: out<=1;
   2180: out<=1;
   2181: out<=1;
   2182: out<=0;
   2183: out<=0;
   2184: out<=0;
   2185: out<=0;
   2186: out<=0;
   2187: out<=0;
   2188: out<=1;
   2189: out<=0;
   2190: out<=0;
   2191: out<=1;
   2192: out<=0;
   2193: out<=1;
   2194: out<=0;
   2195: out<=1;
   2196: out<=1;
   2197: out<=1;
   2198: out<=0;
   2199: out<=0;
   2200: out<=0;
   2201: out<=0;
   2202: out<=0;
   2203: out<=0;
   2204: out<=1;
   2205: out<=0;
   2206: out<=0;
   2207: out<=1;
   2208: out<=0;
   2209: out<=1;
   2210: out<=0;
   2211: out<=1;
   2212: out<=1;
   2213: out<=1;
   2214: out<=0;
   2215: out<=0;
   2216: out<=0;
   2217: out<=0;
   2218: out<=0;
   2219: out<=0;
   2220: out<=1;
   2221: out<=0;
   2222: out<=0;
   2223: out<=1;
   2224: out<=0;
   2225: out<=1;
   2226: out<=0;
   2227: out<=1;
   2228: out<=1;
   2229: out<=1;
   2230: out<=0;
   2231: out<=0;
   2232: out<=0;
   2233: out<=0;
   2234: out<=0;
   2235: out<=0;
   2236: out<=1;
   2237: out<=0;
   2238: out<=0;
   2239: out<=1;
   2240: out<=1;
   2241: out<=0;
   2242: out<=1;
   2243: out<=0;
   2244: out<=0;
   2245: out<=0;
   2246: out<=1;
   2247: out<=1;
   2248: out<=1;
   2249: out<=1;
   2250: out<=1;
   2251: out<=1;
   2252: out<=0;
   2253: out<=1;
   2254: out<=1;
   2255: out<=0;
   2256: out<=0;
   2257: out<=1;
   2258: out<=0;
   2259: out<=1;
   2260: out<=1;
   2261: out<=1;
   2262: out<=0;
   2263: out<=0;
   2264: out<=0;
   2265: out<=0;
   2266: out<=0;
   2267: out<=0;
   2268: out<=1;
   2269: out<=0;
   2270: out<=0;
   2271: out<=1;
   2272: out<=0;
   2273: out<=1;
   2274: out<=0;
   2275: out<=1;
   2276: out<=1;
   2277: out<=1;
   2278: out<=0;
   2279: out<=0;
   2280: out<=0;
   2281: out<=0;
   2282: out<=0;
   2283: out<=0;
   2284: out<=1;
   2285: out<=0;
   2286: out<=0;
   2287: out<=1;
   2288: out<=1;
   2289: out<=0;
   2290: out<=1;
   2291: out<=0;
   2292: out<=0;
   2293: out<=0;
   2294: out<=1;
   2295: out<=1;
   2296: out<=1;
   2297: out<=1;
   2298: out<=1;
   2299: out<=1;
   2300: out<=0;
   2301: out<=1;
   2302: out<=1;
   2303: out<=0;
   2304: out<=1;
   2305: out<=1;
   2306: out<=0;
   2307: out<=0;
   2308: out<=1;
   2309: out<=0;
   2310: out<=1;
   2311: out<=0;
   2312: out<=0;
   2313: out<=1;
   2314: out<=1;
   2315: out<=0;
   2316: out<=0;
   2317: out<=0;
   2318: out<=0;
   2319: out<=0;
   2320: out<=1;
   2321: out<=1;
   2322: out<=0;
   2323: out<=0;
   2324: out<=1;
   2325: out<=0;
   2326: out<=1;
   2327: out<=0;
   2328: out<=0;
   2329: out<=1;
   2330: out<=1;
   2331: out<=0;
   2332: out<=0;
   2333: out<=0;
   2334: out<=0;
   2335: out<=0;
   2336: out<=0;
   2337: out<=0;
   2338: out<=1;
   2339: out<=1;
   2340: out<=0;
   2341: out<=1;
   2342: out<=0;
   2343: out<=1;
   2344: out<=1;
   2345: out<=0;
   2346: out<=0;
   2347: out<=1;
   2348: out<=1;
   2349: out<=1;
   2350: out<=1;
   2351: out<=1;
   2352: out<=0;
   2353: out<=0;
   2354: out<=1;
   2355: out<=1;
   2356: out<=0;
   2357: out<=1;
   2358: out<=0;
   2359: out<=1;
   2360: out<=1;
   2361: out<=0;
   2362: out<=0;
   2363: out<=1;
   2364: out<=1;
   2365: out<=1;
   2366: out<=1;
   2367: out<=1;
   2368: out<=0;
   2369: out<=0;
   2370: out<=1;
   2371: out<=1;
   2372: out<=0;
   2373: out<=1;
   2374: out<=0;
   2375: out<=1;
   2376: out<=1;
   2377: out<=0;
   2378: out<=0;
   2379: out<=1;
   2380: out<=1;
   2381: out<=1;
   2382: out<=1;
   2383: out<=1;
   2384: out<=1;
   2385: out<=1;
   2386: out<=0;
   2387: out<=0;
   2388: out<=1;
   2389: out<=0;
   2390: out<=1;
   2391: out<=0;
   2392: out<=0;
   2393: out<=1;
   2394: out<=1;
   2395: out<=0;
   2396: out<=0;
   2397: out<=0;
   2398: out<=0;
   2399: out<=0;
   2400: out<=0;
   2401: out<=0;
   2402: out<=1;
   2403: out<=1;
   2404: out<=0;
   2405: out<=1;
   2406: out<=0;
   2407: out<=1;
   2408: out<=1;
   2409: out<=0;
   2410: out<=0;
   2411: out<=1;
   2412: out<=1;
   2413: out<=1;
   2414: out<=1;
   2415: out<=1;
   2416: out<=1;
   2417: out<=1;
   2418: out<=0;
   2419: out<=0;
   2420: out<=1;
   2421: out<=0;
   2422: out<=1;
   2423: out<=0;
   2424: out<=0;
   2425: out<=1;
   2426: out<=1;
   2427: out<=0;
   2428: out<=0;
   2429: out<=0;
   2430: out<=0;
   2431: out<=0;
   2432: out<=1;
   2433: out<=1;
   2434: out<=0;
   2435: out<=0;
   2436: out<=1;
   2437: out<=0;
   2438: out<=1;
   2439: out<=0;
   2440: out<=0;
   2441: out<=1;
   2442: out<=1;
   2443: out<=0;
   2444: out<=0;
   2445: out<=0;
   2446: out<=0;
   2447: out<=0;
   2448: out<=0;
   2449: out<=0;
   2450: out<=1;
   2451: out<=1;
   2452: out<=0;
   2453: out<=1;
   2454: out<=0;
   2455: out<=1;
   2456: out<=1;
   2457: out<=0;
   2458: out<=0;
   2459: out<=1;
   2460: out<=1;
   2461: out<=1;
   2462: out<=1;
   2463: out<=1;
   2464: out<=0;
   2465: out<=0;
   2466: out<=1;
   2467: out<=1;
   2468: out<=0;
   2469: out<=1;
   2470: out<=0;
   2471: out<=1;
   2472: out<=1;
   2473: out<=0;
   2474: out<=0;
   2475: out<=1;
   2476: out<=1;
   2477: out<=1;
   2478: out<=1;
   2479: out<=1;
   2480: out<=1;
   2481: out<=1;
   2482: out<=0;
   2483: out<=0;
   2484: out<=1;
   2485: out<=0;
   2486: out<=1;
   2487: out<=0;
   2488: out<=0;
   2489: out<=1;
   2490: out<=1;
   2491: out<=0;
   2492: out<=0;
   2493: out<=0;
   2494: out<=0;
   2495: out<=0;
   2496: out<=0;
   2497: out<=0;
   2498: out<=1;
   2499: out<=1;
   2500: out<=0;
   2501: out<=1;
   2502: out<=0;
   2503: out<=1;
   2504: out<=1;
   2505: out<=0;
   2506: out<=0;
   2507: out<=1;
   2508: out<=1;
   2509: out<=1;
   2510: out<=1;
   2511: out<=1;
   2512: out<=0;
   2513: out<=0;
   2514: out<=1;
   2515: out<=1;
   2516: out<=0;
   2517: out<=1;
   2518: out<=0;
   2519: out<=1;
   2520: out<=1;
   2521: out<=0;
   2522: out<=0;
   2523: out<=1;
   2524: out<=1;
   2525: out<=1;
   2526: out<=1;
   2527: out<=1;
   2528: out<=0;
   2529: out<=0;
   2530: out<=1;
   2531: out<=1;
   2532: out<=0;
   2533: out<=1;
   2534: out<=0;
   2535: out<=1;
   2536: out<=1;
   2537: out<=0;
   2538: out<=0;
   2539: out<=1;
   2540: out<=1;
   2541: out<=1;
   2542: out<=1;
   2543: out<=1;
   2544: out<=0;
   2545: out<=0;
   2546: out<=1;
   2547: out<=1;
   2548: out<=0;
   2549: out<=1;
   2550: out<=0;
   2551: out<=1;
   2552: out<=1;
   2553: out<=0;
   2554: out<=0;
   2555: out<=1;
   2556: out<=1;
   2557: out<=1;
   2558: out<=1;
   2559: out<=1;
   2560: out<=0;
   2561: out<=0;
   2562: out<=0;
   2563: out<=0;
   2564: out<=0;
   2565: out<=1;
   2566: out<=1;
   2567: out<=0;
   2568: out<=0;
   2569: out<=1;
   2570: out<=0;
   2571: out<=1;
   2572: out<=0;
   2573: out<=0;
   2574: out<=1;
   2575: out<=1;
   2576: out<=0;
   2577: out<=0;
   2578: out<=0;
   2579: out<=0;
   2580: out<=0;
   2581: out<=1;
   2582: out<=1;
   2583: out<=0;
   2584: out<=0;
   2585: out<=1;
   2586: out<=0;
   2587: out<=1;
   2588: out<=0;
   2589: out<=0;
   2590: out<=1;
   2591: out<=1;
   2592: out<=0;
   2593: out<=0;
   2594: out<=0;
   2595: out<=0;
   2596: out<=0;
   2597: out<=1;
   2598: out<=1;
   2599: out<=0;
   2600: out<=0;
   2601: out<=1;
   2602: out<=0;
   2603: out<=1;
   2604: out<=0;
   2605: out<=0;
   2606: out<=1;
   2607: out<=1;
   2608: out<=0;
   2609: out<=0;
   2610: out<=0;
   2611: out<=0;
   2612: out<=0;
   2613: out<=1;
   2614: out<=1;
   2615: out<=0;
   2616: out<=0;
   2617: out<=1;
   2618: out<=0;
   2619: out<=1;
   2620: out<=0;
   2621: out<=0;
   2622: out<=1;
   2623: out<=1;
   2624: out<=1;
   2625: out<=1;
   2626: out<=1;
   2627: out<=1;
   2628: out<=1;
   2629: out<=0;
   2630: out<=0;
   2631: out<=1;
   2632: out<=1;
   2633: out<=0;
   2634: out<=1;
   2635: out<=0;
   2636: out<=1;
   2637: out<=1;
   2638: out<=0;
   2639: out<=0;
   2640: out<=0;
   2641: out<=0;
   2642: out<=0;
   2643: out<=0;
   2644: out<=0;
   2645: out<=1;
   2646: out<=1;
   2647: out<=0;
   2648: out<=0;
   2649: out<=1;
   2650: out<=0;
   2651: out<=1;
   2652: out<=0;
   2653: out<=0;
   2654: out<=1;
   2655: out<=1;
   2656: out<=0;
   2657: out<=0;
   2658: out<=0;
   2659: out<=0;
   2660: out<=0;
   2661: out<=1;
   2662: out<=1;
   2663: out<=0;
   2664: out<=0;
   2665: out<=1;
   2666: out<=0;
   2667: out<=1;
   2668: out<=0;
   2669: out<=0;
   2670: out<=1;
   2671: out<=1;
   2672: out<=1;
   2673: out<=1;
   2674: out<=1;
   2675: out<=1;
   2676: out<=1;
   2677: out<=0;
   2678: out<=0;
   2679: out<=1;
   2680: out<=1;
   2681: out<=0;
   2682: out<=1;
   2683: out<=0;
   2684: out<=1;
   2685: out<=1;
   2686: out<=0;
   2687: out<=0;
   2688: out<=0;
   2689: out<=0;
   2690: out<=0;
   2691: out<=0;
   2692: out<=0;
   2693: out<=1;
   2694: out<=1;
   2695: out<=0;
   2696: out<=0;
   2697: out<=1;
   2698: out<=0;
   2699: out<=1;
   2700: out<=0;
   2701: out<=0;
   2702: out<=1;
   2703: out<=1;
   2704: out<=1;
   2705: out<=1;
   2706: out<=1;
   2707: out<=1;
   2708: out<=1;
   2709: out<=0;
   2710: out<=0;
   2711: out<=1;
   2712: out<=1;
   2713: out<=0;
   2714: out<=1;
   2715: out<=0;
   2716: out<=1;
   2717: out<=1;
   2718: out<=0;
   2719: out<=0;
   2720: out<=0;
   2721: out<=0;
   2722: out<=0;
   2723: out<=0;
   2724: out<=0;
   2725: out<=1;
   2726: out<=1;
   2727: out<=0;
   2728: out<=0;
   2729: out<=1;
   2730: out<=0;
   2731: out<=1;
   2732: out<=0;
   2733: out<=0;
   2734: out<=1;
   2735: out<=1;
   2736: out<=1;
   2737: out<=1;
   2738: out<=1;
   2739: out<=1;
   2740: out<=1;
   2741: out<=0;
   2742: out<=0;
   2743: out<=1;
   2744: out<=1;
   2745: out<=0;
   2746: out<=1;
   2747: out<=0;
   2748: out<=1;
   2749: out<=1;
   2750: out<=0;
   2751: out<=0;
   2752: out<=1;
   2753: out<=1;
   2754: out<=1;
   2755: out<=1;
   2756: out<=1;
   2757: out<=0;
   2758: out<=0;
   2759: out<=1;
   2760: out<=1;
   2761: out<=0;
   2762: out<=1;
   2763: out<=0;
   2764: out<=1;
   2765: out<=1;
   2766: out<=0;
   2767: out<=0;
   2768: out<=1;
   2769: out<=1;
   2770: out<=1;
   2771: out<=1;
   2772: out<=1;
   2773: out<=0;
   2774: out<=0;
   2775: out<=1;
   2776: out<=1;
   2777: out<=0;
   2778: out<=1;
   2779: out<=0;
   2780: out<=1;
   2781: out<=1;
   2782: out<=0;
   2783: out<=0;
   2784: out<=0;
   2785: out<=0;
   2786: out<=0;
   2787: out<=0;
   2788: out<=0;
   2789: out<=1;
   2790: out<=1;
   2791: out<=0;
   2792: out<=0;
   2793: out<=1;
   2794: out<=0;
   2795: out<=1;
   2796: out<=0;
   2797: out<=0;
   2798: out<=1;
   2799: out<=1;
   2800: out<=0;
   2801: out<=0;
   2802: out<=0;
   2803: out<=0;
   2804: out<=0;
   2805: out<=1;
   2806: out<=1;
   2807: out<=0;
   2808: out<=0;
   2809: out<=1;
   2810: out<=0;
   2811: out<=1;
   2812: out<=0;
   2813: out<=0;
   2814: out<=1;
   2815: out<=1;
   2816: out<=1;
   2817: out<=0;
   2818: out<=0;
   2819: out<=1;
   2820: out<=0;
   2821: out<=0;
   2822: out<=0;
   2823: out<=0;
   2824: out<=0;
   2825: out<=0;
   2826: out<=1;
   2827: out<=1;
   2828: out<=1;
   2829: out<=0;
   2830: out<=1;
   2831: out<=0;
   2832: out<=0;
   2833: out<=1;
   2834: out<=1;
   2835: out<=0;
   2836: out<=1;
   2837: out<=1;
   2838: out<=1;
   2839: out<=1;
   2840: out<=1;
   2841: out<=1;
   2842: out<=0;
   2843: out<=0;
   2844: out<=0;
   2845: out<=1;
   2846: out<=0;
   2847: out<=1;
   2848: out<=0;
   2849: out<=1;
   2850: out<=1;
   2851: out<=0;
   2852: out<=1;
   2853: out<=1;
   2854: out<=1;
   2855: out<=1;
   2856: out<=1;
   2857: out<=1;
   2858: out<=0;
   2859: out<=0;
   2860: out<=0;
   2861: out<=1;
   2862: out<=0;
   2863: out<=1;
   2864: out<=1;
   2865: out<=0;
   2866: out<=0;
   2867: out<=1;
   2868: out<=0;
   2869: out<=0;
   2870: out<=0;
   2871: out<=0;
   2872: out<=0;
   2873: out<=0;
   2874: out<=1;
   2875: out<=1;
   2876: out<=1;
   2877: out<=0;
   2878: out<=1;
   2879: out<=0;
   2880: out<=0;
   2881: out<=1;
   2882: out<=1;
   2883: out<=0;
   2884: out<=1;
   2885: out<=1;
   2886: out<=1;
   2887: out<=1;
   2888: out<=1;
   2889: out<=1;
   2890: out<=0;
   2891: out<=0;
   2892: out<=0;
   2893: out<=1;
   2894: out<=0;
   2895: out<=1;
   2896: out<=0;
   2897: out<=1;
   2898: out<=1;
   2899: out<=0;
   2900: out<=1;
   2901: out<=1;
   2902: out<=1;
   2903: out<=1;
   2904: out<=1;
   2905: out<=1;
   2906: out<=0;
   2907: out<=0;
   2908: out<=0;
   2909: out<=1;
   2910: out<=0;
   2911: out<=1;
   2912: out<=0;
   2913: out<=1;
   2914: out<=1;
   2915: out<=0;
   2916: out<=1;
   2917: out<=1;
   2918: out<=1;
   2919: out<=1;
   2920: out<=1;
   2921: out<=1;
   2922: out<=0;
   2923: out<=0;
   2924: out<=0;
   2925: out<=1;
   2926: out<=0;
   2927: out<=1;
   2928: out<=0;
   2929: out<=1;
   2930: out<=1;
   2931: out<=0;
   2932: out<=1;
   2933: out<=1;
   2934: out<=1;
   2935: out<=1;
   2936: out<=1;
   2937: out<=1;
   2938: out<=0;
   2939: out<=0;
   2940: out<=0;
   2941: out<=1;
   2942: out<=0;
   2943: out<=1;
   2944: out<=1;
   2945: out<=0;
   2946: out<=0;
   2947: out<=1;
   2948: out<=0;
   2949: out<=0;
   2950: out<=0;
   2951: out<=0;
   2952: out<=0;
   2953: out<=0;
   2954: out<=1;
   2955: out<=1;
   2956: out<=1;
   2957: out<=0;
   2958: out<=1;
   2959: out<=0;
   2960: out<=1;
   2961: out<=0;
   2962: out<=0;
   2963: out<=1;
   2964: out<=0;
   2965: out<=0;
   2966: out<=0;
   2967: out<=0;
   2968: out<=0;
   2969: out<=0;
   2970: out<=1;
   2971: out<=1;
   2972: out<=1;
   2973: out<=0;
   2974: out<=1;
   2975: out<=0;
   2976: out<=0;
   2977: out<=1;
   2978: out<=1;
   2979: out<=0;
   2980: out<=1;
   2981: out<=1;
   2982: out<=1;
   2983: out<=1;
   2984: out<=1;
   2985: out<=1;
   2986: out<=0;
   2987: out<=0;
   2988: out<=0;
   2989: out<=1;
   2990: out<=0;
   2991: out<=1;
   2992: out<=0;
   2993: out<=1;
   2994: out<=1;
   2995: out<=0;
   2996: out<=1;
   2997: out<=1;
   2998: out<=1;
   2999: out<=1;
   3000: out<=1;
   3001: out<=1;
   3002: out<=0;
   3003: out<=0;
   3004: out<=0;
   3005: out<=1;
   3006: out<=0;
   3007: out<=1;
   3008: out<=0;
   3009: out<=1;
   3010: out<=1;
   3011: out<=0;
   3012: out<=1;
   3013: out<=1;
   3014: out<=1;
   3015: out<=1;
   3016: out<=1;
   3017: out<=1;
   3018: out<=0;
   3019: out<=0;
   3020: out<=0;
   3021: out<=1;
   3022: out<=0;
   3023: out<=1;
   3024: out<=1;
   3025: out<=0;
   3026: out<=0;
   3027: out<=1;
   3028: out<=0;
   3029: out<=0;
   3030: out<=0;
   3031: out<=0;
   3032: out<=0;
   3033: out<=0;
   3034: out<=1;
   3035: out<=1;
   3036: out<=1;
   3037: out<=0;
   3038: out<=1;
   3039: out<=0;
   3040: out<=0;
   3041: out<=1;
   3042: out<=1;
   3043: out<=0;
   3044: out<=1;
   3045: out<=1;
   3046: out<=1;
   3047: out<=1;
   3048: out<=1;
   3049: out<=1;
   3050: out<=0;
   3051: out<=0;
   3052: out<=0;
   3053: out<=1;
   3054: out<=0;
   3055: out<=1;
   3056: out<=1;
   3057: out<=0;
   3058: out<=0;
   3059: out<=1;
   3060: out<=0;
   3061: out<=0;
   3062: out<=0;
   3063: out<=0;
   3064: out<=0;
   3065: out<=0;
   3066: out<=1;
   3067: out<=1;
   3068: out<=1;
   3069: out<=0;
   3070: out<=1;
   3071: out<=0;
   3072: out<=0;
   3073: out<=0;
   3074: out<=1;
   3075: out<=1;
   3076: out<=1;
   3077: out<=0;
   3078: out<=1;
   3079: out<=0;
   3080: out<=0;
   3081: out<=1;
   3082: out<=1;
   3083: out<=0;
   3084: out<=1;
   3085: out<=1;
   3086: out<=1;
   3087: out<=1;
   3088: out<=1;
   3089: out<=1;
   3090: out<=0;
   3091: out<=0;
   3092: out<=0;
   3093: out<=1;
   3094: out<=0;
   3095: out<=1;
   3096: out<=1;
   3097: out<=0;
   3098: out<=0;
   3099: out<=1;
   3100: out<=0;
   3101: out<=0;
   3102: out<=0;
   3103: out<=0;
   3104: out<=0;
   3105: out<=0;
   3106: out<=1;
   3107: out<=1;
   3108: out<=1;
   3109: out<=0;
   3110: out<=1;
   3111: out<=0;
   3112: out<=0;
   3113: out<=1;
   3114: out<=1;
   3115: out<=0;
   3116: out<=1;
   3117: out<=1;
   3118: out<=1;
   3119: out<=1;
   3120: out<=1;
   3121: out<=1;
   3122: out<=0;
   3123: out<=0;
   3124: out<=0;
   3125: out<=1;
   3126: out<=0;
   3127: out<=1;
   3128: out<=1;
   3129: out<=0;
   3130: out<=0;
   3131: out<=1;
   3132: out<=0;
   3133: out<=0;
   3134: out<=0;
   3135: out<=0;
   3136: out<=1;
   3137: out<=1;
   3138: out<=0;
   3139: out<=0;
   3140: out<=0;
   3141: out<=1;
   3142: out<=0;
   3143: out<=1;
   3144: out<=1;
   3145: out<=0;
   3146: out<=0;
   3147: out<=1;
   3148: out<=0;
   3149: out<=0;
   3150: out<=0;
   3151: out<=0;
   3152: out<=1;
   3153: out<=1;
   3154: out<=0;
   3155: out<=0;
   3156: out<=0;
   3157: out<=1;
   3158: out<=0;
   3159: out<=1;
   3160: out<=1;
   3161: out<=0;
   3162: out<=0;
   3163: out<=1;
   3164: out<=0;
   3165: out<=0;
   3166: out<=0;
   3167: out<=0;
   3168: out<=0;
   3169: out<=0;
   3170: out<=1;
   3171: out<=1;
   3172: out<=1;
   3173: out<=0;
   3174: out<=1;
   3175: out<=0;
   3176: out<=0;
   3177: out<=1;
   3178: out<=1;
   3179: out<=0;
   3180: out<=1;
   3181: out<=1;
   3182: out<=1;
   3183: out<=1;
   3184: out<=0;
   3185: out<=0;
   3186: out<=1;
   3187: out<=1;
   3188: out<=1;
   3189: out<=0;
   3190: out<=1;
   3191: out<=0;
   3192: out<=0;
   3193: out<=1;
   3194: out<=1;
   3195: out<=0;
   3196: out<=1;
   3197: out<=1;
   3198: out<=1;
   3199: out<=1;
   3200: out<=0;
   3201: out<=0;
   3202: out<=1;
   3203: out<=1;
   3204: out<=1;
   3205: out<=0;
   3206: out<=1;
   3207: out<=0;
   3208: out<=0;
   3209: out<=1;
   3210: out<=1;
   3211: out<=0;
   3212: out<=1;
   3213: out<=1;
   3214: out<=1;
   3215: out<=1;
   3216: out<=0;
   3217: out<=0;
   3218: out<=1;
   3219: out<=1;
   3220: out<=1;
   3221: out<=0;
   3222: out<=1;
   3223: out<=0;
   3224: out<=0;
   3225: out<=1;
   3226: out<=1;
   3227: out<=0;
   3228: out<=1;
   3229: out<=1;
   3230: out<=1;
   3231: out<=1;
   3232: out<=0;
   3233: out<=0;
   3234: out<=1;
   3235: out<=1;
   3236: out<=1;
   3237: out<=0;
   3238: out<=1;
   3239: out<=0;
   3240: out<=0;
   3241: out<=1;
   3242: out<=1;
   3243: out<=0;
   3244: out<=1;
   3245: out<=1;
   3246: out<=1;
   3247: out<=1;
   3248: out<=0;
   3249: out<=0;
   3250: out<=1;
   3251: out<=1;
   3252: out<=1;
   3253: out<=0;
   3254: out<=1;
   3255: out<=0;
   3256: out<=0;
   3257: out<=1;
   3258: out<=1;
   3259: out<=0;
   3260: out<=1;
   3261: out<=1;
   3262: out<=1;
   3263: out<=1;
   3264: out<=1;
   3265: out<=1;
   3266: out<=0;
   3267: out<=0;
   3268: out<=0;
   3269: out<=1;
   3270: out<=0;
   3271: out<=1;
   3272: out<=1;
   3273: out<=0;
   3274: out<=0;
   3275: out<=1;
   3276: out<=0;
   3277: out<=0;
   3278: out<=0;
   3279: out<=0;
   3280: out<=0;
   3281: out<=0;
   3282: out<=1;
   3283: out<=1;
   3284: out<=1;
   3285: out<=0;
   3286: out<=1;
   3287: out<=0;
   3288: out<=0;
   3289: out<=1;
   3290: out<=1;
   3291: out<=0;
   3292: out<=1;
   3293: out<=1;
   3294: out<=1;
   3295: out<=1;
   3296: out<=0;
   3297: out<=0;
   3298: out<=1;
   3299: out<=1;
   3300: out<=1;
   3301: out<=0;
   3302: out<=1;
   3303: out<=0;
   3304: out<=0;
   3305: out<=1;
   3306: out<=1;
   3307: out<=0;
   3308: out<=1;
   3309: out<=1;
   3310: out<=1;
   3311: out<=1;
   3312: out<=1;
   3313: out<=1;
   3314: out<=0;
   3315: out<=0;
   3316: out<=0;
   3317: out<=1;
   3318: out<=0;
   3319: out<=1;
   3320: out<=1;
   3321: out<=0;
   3322: out<=0;
   3323: out<=1;
   3324: out<=0;
   3325: out<=0;
   3326: out<=0;
   3327: out<=0;
   3328: out<=0;
   3329: out<=1;
   3330: out<=0;
   3331: out<=1;
   3332: out<=0;
   3333: out<=0;
   3334: out<=1;
   3335: out<=1;
   3336: out<=1;
   3337: out<=1;
   3338: out<=1;
   3339: out<=1;
   3340: out<=1;
   3341: out<=0;
   3342: out<=0;
   3343: out<=1;
   3344: out<=0;
   3345: out<=1;
   3346: out<=0;
   3347: out<=1;
   3348: out<=0;
   3349: out<=0;
   3350: out<=1;
   3351: out<=1;
   3352: out<=1;
   3353: out<=1;
   3354: out<=1;
   3355: out<=1;
   3356: out<=1;
   3357: out<=0;
   3358: out<=0;
   3359: out<=1;
   3360: out<=1;
   3361: out<=0;
   3362: out<=1;
   3363: out<=0;
   3364: out<=1;
   3365: out<=1;
   3366: out<=0;
   3367: out<=0;
   3368: out<=0;
   3369: out<=0;
   3370: out<=0;
   3371: out<=0;
   3372: out<=0;
   3373: out<=1;
   3374: out<=1;
   3375: out<=0;
   3376: out<=1;
   3377: out<=0;
   3378: out<=1;
   3379: out<=0;
   3380: out<=1;
   3381: out<=1;
   3382: out<=0;
   3383: out<=0;
   3384: out<=0;
   3385: out<=0;
   3386: out<=0;
   3387: out<=0;
   3388: out<=0;
   3389: out<=1;
   3390: out<=1;
   3391: out<=0;
   3392: out<=1;
   3393: out<=0;
   3394: out<=1;
   3395: out<=0;
   3396: out<=1;
   3397: out<=1;
   3398: out<=0;
   3399: out<=0;
   3400: out<=0;
   3401: out<=0;
   3402: out<=0;
   3403: out<=0;
   3404: out<=0;
   3405: out<=1;
   3406: out<=1;
   3407: out<=0;
   3408: out<=0;
   3409: out<=1;
   3410: out<=0;
   3411: out<=1;
   3412: out<=0;
   3413: out<=0;
   3414: out<=1;
   3415: out<=1;
   3416: out<=1;
   3417: out<=1;
   3418: out<=1;
   3419: out<=1;
   3420: out<=1;
   3421: out<=0;
   3422: out<=0;
   3423: out<=1;
   3424: out<=1;
   3425: out<=0;
   3426: out<=1;
   3427: out<=0;
   3428: out<=1;
   3429: out<=1;
   3430: out<=0;
   3431: out<=0;
   3432: out<=0;
   3433: out<=0;
   3434: out<=0;
   3435: out<=0;
   3436: out<=0;
   3437: out<=1;
   3438: out<=1;
   3439: out<=0;
   3440: out<=0;
   3441: out<=1;
   3442: out<=0;
   3443: out<=1;
   3444: out<=0;
   3445: out<=0;
   3446: out<=1;
   3447: out<=1;
   3448: out<=1;
   3449: out<=1;
   3450: out<=1;
   3451: out<=1;
   3452: out<=1;
   3453: out<=0;
   3454: out<=0;
   3455: out<=1;
   3456: out<=0;
   3457: out<=1;
   3458: out<=0;
   3459: out<=1;
   3460: out<=0;
   3461: out<=0;
   3462: out<=1;
   3463: out<=1;
   3464: out<=1;
   3465: out<=1;
   3466: out<=1;
   3467: out<=1;
   3468: out<=1;
   3469: out<=0;
   3470: out<=0;
   3471: out<=1;
   3472: out<=1;
   3473: out<=0;
   3474: out<=1;
   3475: out<=0;
   3476: out<=1;
   3477: out<=1;
   3478: out<=0;
   3479: out<=0;
   3480: out<=0;
   3481: out<=0;
   3482: out<=0;
   3483: out<=0;
   3484: out<=0;
   3485: out<=1;
   3486: out<=1;
   3487: out<=0;
   3488: out<=1;
   3489: out<=0;
   3490: out<=1;
   3491: out<=0;
   3492: out<=1;
   3493: out<=1;
   3494: out<=0;
   3495: out<=0;
   3496: out<=0;
   3497: out<=0;
   3498: out<=0;
   3499: out<=0;
   3500: out<=0;
   3501: out<=1;
   3502: out<=1;
   3503: out<=0;
   3504: out<=0;
   3505: out<=1;
   3506: out<=0;
   3507: out<=1;
   3508: out<=0;
   3509: out<=0;
   3510: out<=1;
   3511: out<=1;
   3512: out<=1;
   3513: out<=1;
   3514: out<=1;
   3515: out<=1;
   3516: out<=1;
   3517: out<=0;
   3518: out<=0;
   3519: out<=1;
   3520: out<=1;
   3521: out<=0;
   3522: out<=1;
   3523: out<=0;
   3524: out<=1;
   3525: out<=1;
   3526: out<=0;
   3527: out<=0;
   3528: out<=0;
   3529: out<=0;
   3530: out<=0;
   3531: out<=0;
   3532: out<=0;
   3533: out<=1;
   3534: out<=1;
   3535: out<=0;
   3536: out<=1;
   3537: out<=0;
   3538: out<=1;
   3539: out<=0;
   3540: out<=1;
   3541: out<=1;
   3542: out<=0;
   3543: out<=0;
   3544: out<=0;
   3545: out<=0;
   3546: out<=0;
   3547: out<=0;
   3548: out<=0;
   3549: out<=1;
   3550: out<=1;
   3551: out<=0;
   3552: out<=1;
   3553: out<=0;
   3554: out<=1;
   3555: out<=0;
   3556: out<=1;
   3557: out<=1;
   3558: out<=0;
   3559: out<=0;
   3560: out<=0;
   3561: out<=0;
   3562: out<=0;
   3563: out<=0;
   3564: out<=0;
   3565: out<=1;
   3566: out<=1;
   3567: out<=0;
   3568: out<=1;
   3569: out<=0;
   3570: out<=1;
   3571: out<=0;
   3572: out<=1;
   3573: out<=1;
   3574: out<=0;
   3575: out<=0;
   3576: out<=0;
   3577: out<=0;
   3578: out<=0;
   3579: out<=0;
   3580: out<=0;
   3581: out<=1;
   3582: out<=1;
   3583: out<=0;
   3584: out<=1;
   3585: out<=0;
   3586: out<=0;
   3587: out<=1;
   3588: out<=1;
   3589: out<=1;
   3590: out<=1;
   3591: out<=1;
   3592: out<=1;
   3593: out<=1;
   3594: out<=0;
   3595: out<=0;
   3596: out<=1;
   3597: out<=0;
   3598: out<=1;
   3599: out<=0;
   3600: out<=1;
   3601: out<=0;
   3602: out<=0;
   3603: out<=1;
   3604: out<=1;
   3605: out<=1;
   3606: out<=1;
   3607: out<=1;
   3608: out<=1;
   3609: out<=1;
   3610: out<=0;
   3611: out<=0;
   3612: out<=1;
   3613: out<=0;
   3614: out<=1;
   3615: out<=0;
   3616: out<=1;
   3617: out<=0;
   3618: out<=0;
   3619: out<=1;
   3620: out<=1;
   3621: out<=1;
   3622: out<=1;
   3623: out<=1;
   3624: out<=1;
   3625: out<=1;
   3626: out<=0;
   3627: out<=0;
   3628: out<=1;
   3629: out<=0;
   3630: out<=1;
   3631: out<=0;
   3632: out<=1;
   3633: out<=0;
   3634: out<=0;
   3635: out<=1;
   3636: out<=1;
   3637: out<=1;
   3638: out<=1;
   3639: out<=1;
   3640: out<=1;
   3641: out<=1;
   3642: out<=0;
   3643: out<=0;
   3644: out<=1;
   3645: out<=0;
   3646: out<=1;
   3647: out<=0;
   3648: out<=0;
   3649: out<=1;
   3650: out<=1;
   3651: out<=0;
   3652: out<=0;
   3653: out<=0;
   3654: out<=0;
   3655: out<=0;
   3656: out<=0;
   3657: out<=0;
   3658: out<=1;
   3659: out<=1;
   3660: out<=0;
   3661: out<=1;
   3662: out<=0;
   3663: out<=1;
   3664: out<=1;
   3665: out<=0;
   3666: out<=0;
   3667: out<=1;
   3668: out<=1;
   3669: out<=1;
   3670: out<=1;
   3671: out<=1;
   3672: out<=1;
   3673: out<=1;
   3674: out<=0;
   3675: out<=0;
   3676: out<=1;
   3677: out<=0;
   3678: out<=1;
   3679: out<=0;
   3680: out<=1;
   3681: out<=0;
   3682: out<=0;
   3683: out<=1;
   3684: out<=1;
   3685: out<=1;
   3686: out<=1;
   3687: out<=1;
   3688: out<=1;
   3689: out<=1;
   3690: out<=0;
   3691: out<=0;
   3692: out<=1;
   3693: out<=0;
   3694: out<=1;
   3695: out<=0;
   3696: out<=0;
   3697: out<=1;
   3698: out<=1;
   3699: out<=0;
   3700: out<=0;
   3701: out<=0;
   3702: out<=0;
   3703: out<=0;
   3704: out<=0;
   3705: out<=0;
   3706: out<=1;
   3707: out<=1;
   3708: out<=0;
   3709: out<=1;
   3710: out<=0;
   3711: out<=1;
   3712: out<=1;
   3713: out<=0;
   3714: out<=0;
   3715: out<=1;
   3716: out<=1;
   3717: out<=1;
   3718: out<=1;
   3719: out<=1;
   3720: out<=1;
   3721: out<=1;
   3722: out<=0;
   3723: out<=0;
   3724: out<=1;
   3725: out<=0;
   3726: out<=1;
   3727: out<=0;
   3728: out<=0;
   3729: out<=1;
   3730: out<=1;
   3731: out<=0;
   3732: out<=0;
   3733: out<=0;
   3734: out<=0;
   3735: out<=0;
   3736: out<=0;
   3737: out<=0;
   3738: out<=1;
   3739: out<=1;
   3740: out<=0;
   3741: out<=1;
   3742: out<=0;
   3743: out<=1;
   3744: out<=1;
   3745: out<=0;
   3746: out<=0;
   3747: out<=1;
   3748: out<=1;
   3749: out<=1;
   3750: out<=1;
   3751: out<=1;
   3752: out<=1;
   3753: out<=1;
   3754: out<=0;
   3755: out<=0;
   3756: out<=1;
   3757: out<=0;
   3758: out<=1;
   3759: out<=0;
   3760: out<=0;
   3761: out<=1;
   3762: out<=1;
   3763: out<=0;
   3764: out<=0;
   3765: out<=0;
   3766: out<=0;
   3767: out<=0;
   3768: out<=0;
   3769: out<=0;
   3770: out<=1;
   3771: out<=1;
   3772: out<=0;
   3773: out<=1;
   3774: out<=0;
   3775: out<=1;
   3776: out<=0;
   3777: out<=1;
   3778: out<=1;
   3779: out<=0;
   3780: out<=0;
   3781: out<=0;
   3782: out<=0;
   3783: out<=0;
   3784: out<=0;
   3785: out<=0;
   3786: out<=1;
   3787: out<=1;
   3788: out<=0;
   3789: out<=1;
   3790: out<=0;
   3791: out<=1;
   3792: out<=0;
   3793: out<=1;
   3794: out<=1;
   3795: out<=0;
   3796: out<=0;
   3797: out<=0;
   3798: out<=0;
   3799: out<=0;
   3800: out<=0;
   3801: out<=0;
   3802: out<=1;
   3803: out<=1;
   3804: out<=0;
   3805: out<=1;
   3806: out<=0;
   3807: out<=1;
   3808: out<=1;
   3809: out<=0;
   3810: out<=0;
   3811: out<=1;
   3812: out<=1;
   3813: out<=1;
   3814: out<=1;
   3815: out<=1;
   3816: out<=1;
   3817: out<=1;
   3818: out<=0;
   3819: out<=0;
   3820: out<=1;
   3821: out<=0;
   3822: out<=1;
   3823: out<=0;
   3824: out<=1;
   3825: out<=0;
   3826: out<=0;
   3827: out<=1;
   3828: out<=1;
   3829: out<=1;
   3830: out<=1;
   3831: out<=1;
   3832: out<=1;
   3833: out<=1;
   3834: out<=0;
   3835: out<=0;
   3836: out<=1;
   3837: out<=0;
   3838: out<=1;
   3839: out<=0;
   3840: out<=1;
   3841: out<=1;
   3842: out<=1;
   3843: out<=1;
   3844: out<=0;
   3845: out<=1;
   3846: out<=1;
   3847: out<=0;
   3848: out<=0;
   3849: out<=1;
   3850: out<=0;
   3851: out<=1;
   3852: out<=1;
   3853: out<=1;
   3854: out<=0;
   3855: out<=0;
   3856: out<=0;
   3857: out<=0;
   3858: out<=0;
   3859: out<=0;
   3860: out<=1;
   3861: out<=0;
   3862: out<=0;
   3863: out<=1;
   3864: out<=1;
   3865: out<=0;
   3866: out<=1;
   3867: out<=0;
   3868: out<=0;
   3869: out<=0;
   3870: out<=1;
   3871: out<=1;
   3872: out<=0;
   3873: out<=0;
   3874: out<=0;
   3875: out<=0;
   3876: out<=1;
   3877: out<=0;
   3878: out<=0;
   3879: out<=1;
   3880: out<=1;
   3881: out<=0;
   3882: out<=1;
   3883: out<=0;
   3884: out<=0;
   3885: out<=0;
   3886: out<=1;
   3887: out<=1;
   3888: out<=1;
   3889: out<=1;
   3890: out<=1;
   3891: out<=1;
   3892: out<=0;
   3893: out<=1;
   3894: out<=1;
   3895: out<=0;
   3896: out<=0;
   3897: out<=1;
   3898: out<=0;
   3899: out<=1;
   3900: out<=1;
   3901: out<=1;
   3902: out<=0;
   3903: out<=0;
   3904: out<=0;
   3905: out<=0;
   3906: out<=0;
   3907: out<=0;
   3908: out<=1;
   3909: out<=0;
   3910: out<=0;
   3911: out<=1;
   3912: out<=1;
   3913: out<=0;
   3914: out<=1;
   3915: out<=0;
   3916: out<=0;
   3917: out<=0;
   3918: out<=1;
   3919: out<=1;
   3920: out<=0;
   3921: out<=0;
   3922: out<=0;
   3923: out<=0;
   3924: out<=1;
   3925: out<=0;
   3926: out<=0;
   3927: out<=1;
   3928: out<=1;
   3929: out<=0;
   3930: out<=1;
   3931: out<=0;
   3932: out<=0;
   3933: out<=0;
   3934: out<=1;
   3935: out<=1;
   3936: out<=0;
   3937: out<=0;
   3938: out<=0;
   3939: out<=0;
   3940: out<=1;
   3941: out<=0;
   3942: out<=0;
   3943: out<=1;
   3944: out<=1;
   3945: out<=0;
   3946: out<=1;
   3947: out<=0;
   3948: out<=0;
   3949: out<=0;
   3950: out<=1;
   3951: out<=1;
   3952: out<=0;
   3953: out<=0;
   3954: out<=0;
   3955: out<=0;
   3956: out<=1;
   3957: out<=0;
   3958: out<=0;
   3959: out<=1;
   3960: out<=1;
   3961: out<=0;
   3962: out<=1;
   3963: out<=0;
   3964: out<=0;
   3965: out<=0;
   3966: out<=1;
   3967: out<=1;
   3968: out<=1;
   3969: out<=1;
   3970: out<=1;
   3971: out<=1;
   3972: out<=0;
   3973: out<=1;
   3974: out<=1;
   3975: out<=0;
   3976: out<=0;
   3977: out<=1;
   3978: out<=0;
   3979: out<=1;
   3980: out<=1;
   3981: out<=1;
   3982: out<=0;
   3983: out<=0;
   3984: out<=1;
   3985: out<=1;
   3986: out<=1;
   3987: out<=1;
   3988: out<=0;
   3989: out<=1;
   3990: out<=1;
   3991: out<=0;
   3992: out<=0;
   3993: out<=1;
   3994: out<=0;
   3995: out<=1;
   3996: out<=1;
   3997: out<=1;
   3998: out<=0;
   3999: out<=0;
   4000: out<=0;
   4001: out<=0;
   4002: out<=0;
   4003: out<=0;
   4004: out<=1;
   4005: out<=0;
   4006: out<=0;
   4007: out<=1;
   4008: out<=1;
   4009: out<=0;
   4010: out<=1;
   4011: out<=0;
   4012: out<=0;
   4013: out<=0;
   4014: out<=1;
   4015: out<=1;
   4016: out<=0;
   4017: out<=0;
   4018: out<=0;
   4019: out<=0;
   4020: out<=1;
   4021: out<=0;
   4022: out<=0;
   4023: out<=1;
   4024: out<=1;
   4025: out<=0;
   4026: out<=1;
   4027: out<=0;
   4028: out<=0;
   4029: out<=0;
   4030: out<=1;
   4031: out<=1;
   4032: out<=0;
   4033: out<=0;
   4034: out<=0;
   4035: out<=0;
   4036: out<=1;
   4037: out<=0;
   4038: out<=0;
   4039: out<=1;
   4040: out<=1;
   4041: out<=0;
   4042: out<=1;
   4043: out<=0;
   4044: out<=0;
   4045: out<=0;
   4046: out<=1;
   4047: out<=1;
   4048: out<=1;
   4049: out<=1;
   4050: out<=1;
   4051: out<=1;
   4052: out<=0;
   4053: out<=1;
   4054: out<=1;
   4055: out<=0;
   4056: out<=0;
   4057: out<=1;
   4058: out<=0;
   4059: out<=1;
   4060: out<=1;
   4061: out<=1;
   4062: out<=0;
   4063: out<=0;
   4064: out<=0;
   4065: out<=0;
   4066: out<=0;
   4067: out<=0;
   4068: out<=1;
   4069: out<=0;
   4070: out<=0;
   4071: out<=1;
   4072: out<=1;
   4073: out<=0;
   4074: out<=1;
   4075: out<=0;
   4076: out<=0;
   4077: out<=0;
   4078: out<=1;
   4079: out<=1;
   4080: out<=1;
   4081: out<=1;
   4082: out<=1;
   4083: out<=1;
   4084: out<=0;
   4085: out<=1;
   4086: out<=1;
   4087: out<=0;
   4088: out<=0;
   4089: out<=1;
   4090: out<=0;
   4091: out<=1;
   4092: out<=1;
   4093: out<=1;
   4094: out<=0;
   4095: out<=0;
   4096: out<=0;
   4097: out<=1;
   4098: out<=1;
   4099: out<=0;
   4100: out<=1;
   4101: out<=1;
   4102: out<=1;
   4103: out<=1;
   4104: out<=0;
   4105: out<=0;
   4106: out<=1;
   4107: out<=1;
   4108: out<=1;
   4109: out<=0;
   4110: out<=1;
   4111: out<=0;
   4112: out<=0;
   4113: out<=1;
   4114: out<=1;
   4115: out<=0;
   4116: out<=1;
   4117: out<=1;
   4118: out<=1;
   4119: out<=1;
   4120: out<=0;
   4121: out<=0;
   4122: out<=1;
   4123: out<=1;
   4124: out<=1;
   4125: out<=0;
   4126: out<=1;
   4127: out<=0;
   4128: out<=1;
   4129: out<=0;
   4130: out<=0;
   4131: out<=1;
   4132: out<=0;
   4133: out<=0;
   4134: out<=0;
   4135: out<=0;
   4136: out<=1;
   4137: out<=1;
   4138: out<=0;
   4139: out<=0;
   4140: out<=0;
   4141: out<=1;
   4142: out<=0;
   4143: out<=1;
   4144: out<=1;
   4145: out<=0;
   4146: out<=0;
   4147: out<=1;
   4148: out<=0;
   4149: out<=0;
   4150: out<=0;
   4151: out<=0;
   4152: out<=1;
   4153: out<=1;
   4154: out<=0;
   4155: out<=0;
   4156: out<=0;
   4157: out<=1;
   4158: out<=0;
   4159: out<=1;
   4160: out<=0;
   4161: out<=1;
   4162: out<=1;
   4163: out<=0;
   4164: out<=1;
   4165: out<=1;
   4166: out<=1;
   4167: out<=1;
   4168: out<=0;
   4169: out<=0;
   4170: out<=1;
   4171: out<=1;
   4172: out<=1;
   4173: out<=0;
   4174: out<=1;
   4175: out<=0;
   4176: out<=1;
   4177: out<=0;
   4178: out<=0;
   4179: out<=1;
   4180: out<=0;
   4181: out<=0;
   4182: out<=0;
   4183: out<=0;
   4184: out<=1;
   4185: out<=1;
   4186: out<=0;
   4187: out<=0;
   4188: out<=0;
   4189: out<=1;
   4190: out<=0;
   4191: out<=1;
   4192: out<=0;
   4193: out<=1;
   4194: out<=1;
   4195: out<=0;
   4196: out<=1;
   4197: out<=1;
   4198: out<=1;
   4199: out<=1;
   4200: out<=0;
   4201: out<=0;
   4202: out<=1;
   4203: out<=1;
   4204: out<=1;
   4205: out<=0;
   4206: out<=1;
   4207: out<=0;
   4208: out<=1;
   4209: out<=0;
   4210: out<=0;
   4211: out<=1;
   4212: out<=0;
   4213: out<=0;
   4214: out<=0;
   4215: out<=0;
   4216: out<=1;
   4217: out<=1;
   4218: out<=0;
   4219: out<=0;
   4220: out<=0;
   4221: out<=1;
   4222: out<=0;
   4223: out<=1;
   4224: out<=1;
   4225: out<=0;
   4226: out<=0;
   4227: out<=1;
   4228: out<=0;
   4229: out<=0;
   4230: out<=0;
   4231: out<=0;
   4232: out<=1;
   4233: out<=1;
   4234: out<=0;
   4235: out<=0;
   4236: out<=0;
   4237: out<=1;
   4238: out<=0;
   4239: out<=1;
   4240: out<=0;
   4241: out<=1;
   4242: out<=1;
   4243: out<=0;
   4244: out<=1;
   4245: out<=1;
   4246: out<=1;
   4247: out<=1;
   4248: out<=0;
   4249: out<=0;
   4250: out<=1;
   4251: out<=1;
   4252: out<=1;
   4253: out<=0;
   4254: out<=1;
   4255: out<=0;
   4256: out<=0;
   4257: out<=1;
   4258: out<=1;
   4259: out<=0;
   4260: out<=1;
   4261: out<=1;
   4262: out<=1;
   4263: out<=1;
   4264: out<=0;
   4265: out<=0;
   4266: out<=1;
   4267: out<=1;
   4268: out<=1;
   4269: out<=0;
   4270: out<=1;
   4271: out<=0;
   4272: out<=1;
   4273: out<=0;
   4274: out<=0;
   4275: out<=1;
   4276: out<=0;
   4277: out<=0;
   4278: out<=0;
   4279: out<=0;
   4280: out<=1;
   4281: out<=1;
   4282: out<=0;
   4283: out<=0;
   4284: out<=0;
   4285: out<=1;
   4286: out<=0;
   4287: out<=1;
   4288: out<=1;
   4289: out<=0;
   4290: out<=0;
   4291: out<=1;
   4292: out<=0;
   4293: out<=0;
   4294: out<=0;
   4295: out<=0;
   4296: out<=1;
   4297: out<=1;
   4298: out<=0;
   4299: out<=0;
   4300: out<=0;
   4301: out<=1;
   4302: out<=0;
   4303: out<=1;
   4304: out<=1;
   4305: out<=0;
   4306: out<=0;
   4307: out<=1;
   4308: out<=0;
   4309: out<=0;
   4310: out<=0;
   4311: out<=0;
   4312: out<=1;
   4313: out<=1;
   4314: out<=0;
   4315: out<=0;
   4316: out<=0;
   4317: out<=1;
   4318: out<=0;
   4319: out<=1;
   4320: out<=1;
   4321: out<=0;
   4322: out<=0;
   4323: out<=1;
   4324: out<=0;
   4325: out<=0;
   4326: out<=0;
   4327: out<=0;
   4328: out<=1;
   4329: out<=1;
   4330: out<=0;
   4331: out<=0;
   4332: out<=0;
   4333: out<=1;
   4334: out<=0;
   4335: out<=1;
   4336: out<=1;
   4337: out<=0;
   4338: out<=0;
   4339: out<=1;
   4340: out<=0;
   4341: out<=0;
   4342: out<=0;
   4343: out<=0;
   4344: out<=1;
   4345: out<=1;
   4346: out<=0;
   4347: out<=0;
   4348: out<=0;
   4349: out<=1;
   4350: out<=0;
   4351: out<=1;
   4352: out<=0;
   4353: out<=0;
   4354: out<=0;
   4355: out<=0;
   4356: out<=0;
   4357: out<=1;
   4358: out<=1;
   4359: out<=0;
   4360: out<=1;
   4361: out<=0;
   4362: out<=1;
   4363: out<=0;
   4364: out<=1;
   4365: out<=1;
   4366: out<=0;
   4367: out<=0;
   4368: out<=1;
   4369: out<=1;
   4370: out<=1;
   4371: out<=1;
   4372: out<=1;
   4373: out<=0;
   4374: out<=0;
   4375: out<=1;
   4376: out<=0;
   4377: out<=1;
   4378: out<=0;
   4379: out<=1;
   4380: out<=0;
   4381: out<=0;
   4382: out<=1;
   4383: out<=1;
   4384: out<=0;
   4385: out<=0;
   4386: out<=0;
   4387: out<=0;
   4388: out<=0;
   4389: out<=1;
   4390: out<=1;
   4391: out<=0;
   4392: out<=1;
   4393: out<=0;
   4394: out<=1;
   4395: out<=0;
   4396: out<=1;
   4397: out<=1;
   4398: out<=0;
   4399: out<=0;
   4400: out<=1;
   4401: out<=1;
   4402: out<=1;
   4403: out<=1;
   4404: out<=1;
   4405: out<=0;
   4406: out<=0;
   4407: out<=1;
   4408: out<=0;
   4409: out<=1;
   4410: out<=0;
   4411: out<=1;
   4412: out<=0;
   4413: out<=0;
   4414: out<=1;
   4415: out<=1;
   4416: out<=0;
   4417: out<=0;
   4418: out<=0;
   4419: out<=0;
   4420: out<=0;
   4421: out<=1;
   4422: out<=1;
   4423: out<=0;
   4424: out<=1;
   4425: out<=0;
   4426: out<=1;
   4427: out<=0;
   4428: out<=1;
   4429: out<=1;
   4430: out<=0;
   4431: out<=0;
   4432: out<=0;
   4433: out<=0;
   4434: out<=0;
   4435: out<=0;
   4436: out<=0;
   4437: out<=1;
   4438: out<=1;
   4439: out<=0;
   4440: out<=1;
   4441: out<=0;
   4442: out<=1;
   4443: out<=0;
   4444: out<=1;
   4445: out<=1;
   4446: out<=0;
   4447: out<=0;
   4448: out<=1;
   4449: out<=1;
   4450: out<=1;
   4451: out<=1;
   4452: out<=1;
   4453: out<=0;
   4454: out<=0;
   4455: out<=1;
   4456: out<=0;
   4457: out<=1;
   4458: out<=0;
   4459: out<=1;
   4460: out<=0;
   4461: out<=0;
   4462: out<=1;
   4463: out<=1;
   4464: out<=1;
   4465: out<=1;
   4466: out<=1;
   4467: out<=1;
   4468: out<=1;
   4469: out<=0;
   4470: out<=0;
   4471: out<=1;
   4472: out<=0;
   4473: out<=1;
   4474: out<=0;
   4475: out<=1;
   4476: out<=0;
   4477: out<=0;
   4478: out<=1;
   4479: out<=1;
   4480: out<=1;
   4481: out<=1;
   4482: out<=1;
   4483: out<=1;
   4484: out<=1;
   4485: out<=0;
   4486: out<=0;
   4487: out<=1;
   4488: out<=0;
   4489: out<=1;
   4490: out<=0;
   4491: out<=1;
   4492: out<=0;
   4493: out<=0;
   4494: out<=1;
   4495: out<=1;
   4496: out<=1;
   4497: out<=1;
   4498: out<=1;
   4499: out<=1;
   4500: out<=1;
   4501: out<=0;
   4502: out<=0;
   4503: out<=1;
   4504: out<=0;
   4505: out<=1;
   4506: out<=0;
   4507: out<=1;
   4508: out<=0;
   4509: out<=0;
   4510: out<=1;
   4511: out<=1;
   4512: out<=1;
   4513: out<=1;
   4514: out<=1;
   4515: out<=1;
   4516: out<=1;
   4517: out<=0;
   4518: out<=0;
   4519: out<=1;
   4520: out<=0;
   4521: out<=1;
   4522: out<=0;
   4523: out<=1;
   4524: out<=0;
   4525: out<=0;
   4526: out<=1;
   4527: out<=1;
   4528: out<=1;
   4529: out<=1;
   4530: out<=1;
   4531: out<=1;
   4532: out<=1;
   4533: out<=0;
   4534: out<=0;
   4535: out<=1;
   4536: out<=0;
   4537: out<=1;
   4538: out<=0;
   4539: out<=1;
   4540: out<=0;
   4541: out<=0;
   4542: out<=1;
   4543: out<=1;
   4544: out<=1;
   4545: out<=1;
   4546: out<=1;
   4547: out<=1;
   4548: out<=1;
   4549: out<=0;
   4550: out<=0;
   4551: out<=1;
   4552: out<=0;
   4553: out<=1;
   4554: out<=0;
   4555: out<=1;
   4556: out<=0;
   4557: out<=0;
   4558: out<=1;
   4559: out<=1;
   4560: out<=0;
   4561: out<=0;
   4562: out<=0;
   4563: out<=0;
   4564: out<=0;
   4565: out<=1;
   4566: out<=1;
   4567: out<=0;
   4568: out<=1;
   4569: out<=0;
   4570: out<=1;
   4571: out<=0;
   4572: out<=1;
   4573: out<=1;
   4574: out<=0;
   4575: out<=0;
   4576: out<=0;
   4577: out<=0;
   4578: out<=0;
   4579: out<=0;
   4580: out<=0;
   4581: out<=1;
   4582: out<=1;
   4583: out<=0;
   4584: out<=1;
   4585: out<=0;
   4586: out<=1;
   4587: out<=0;
   4588: out<=1;
   4589: out<=1;
   4590: out<=0;
   4591: out<=0;
   4592: out<=1;
   4593: out<=1;
   4594: out<=1;
   4595: out<=1;
   4596: out<=1;
   4597: out<=0;
   4598: out<=0;
   4599: out<=1;
   4600: out<=0;
   4601: out<=1;
   4602: out<=0;
   4603: out<=1;
   4604: out<=0;
   4605: out<=0;
   4606: out<=1;
   4607: out<=1;
   4608: out<=0;
   4609: out<=0;
   4610: out<=1;
   4611: out<=1;
   4612: out<=0;
   4613: out<=1;
   4614: out<=0;
   4615: out<=1;
   4616: out<=0;
   4617: out<=1;
   4618: out<=1;
   4619: out<=0;
   4620: out<=0;
   4621: out<=0;
   4622: out<=0;
   4623: out<=0;
   4624: out<=1;
   4625: out<=1;
   4626: out<=0;
   4627: out<=0;
   4628: out<=1;
   4629: out<=0;
   4630: out<=1;
   4631: out<=0;
   4632: out<=1;
   4633: out<=0;
   4634: out<=0;
   4635: out<=1;
   4636: out<=1;
   4637: out<=1;
   4638: out<=1;
   4639: out<=1;
   4640: out<=1;
   4641: out<=1;
   4642: out<=0;
   4643: out<=0;
   4644: out<=1;
   4645: out<=0;
   4646: out<=1;
   4647: out<=0;
   4648: out<=1;
   4649: out<=0;
   4650: out<=0;
   4651: out<=1;
   4652: out<=1;
   4653: out<=1;
   4654: out<=1;
   4655: out<=1;
   4656: out<=0;
   4657: out<=0;
   4658: out<=1;
   4659: out<=1;
   4660: out<=0;
   4661: out<=1;
   4662: out<=0;
   4663: out<=1;
   4664: out<=0;
   4665: out<=1;
   4666: out<=1;
   4667: out<=0;
   4668: out<=0;
   4669: out<=0;
   4670: out<=0;
   4671: out<=0;
   4672: out<=0;
   4673: out<=0;
   4674: out<=1;
   4675: out<=1;
   4676: out<=0;
   4677: out<=1;
   4678: out<=0;
   4679: out<=1;
   4680: out<=0;
   4681: out<=1;
   4682: out<=1;
   4683: out<=0;
   4684: out<=0;
   4685: out<=0;
   4686: out<=0;
   4687: out<=0;
   4688: out<=0;
   4689: out<=0;
   4690: out<=1;
   4691: out<=1;
   4692: out<=0;
   4693: out<=1;
   4694: out<=0;
   4695: out<=1;
   4696: out<=0;
   4697: out<=1;
   4698: out<=1;
   4699: out<=0;
   4700: out<=0;
   4701: out<=0;
   4702: out<=0;
   4703: out<=0;
   4704: out<=0;
   4705: out<=0;
   4706: out<=1;
   4707: out<=1;
   4708: out<=0;
   4709: out<=1;
   4710: out<=0;
   4711: out<=1;
   4712: out<=0;
   4713: out<=1;
   4714: out<=1;
   4715: out<=0;
   4716: out<=0;
   4717: out<=0;
   4718: out<=0;
   4719: out<=0;
   4720: out<=0;
   4721: out<=0;
   4722: out<=1;
   4723: out<=1;
   4724: out<=0;
   4725: out<=1;
   4726: out<=0;
   4727: out<=1;
   4728: out<=0;
   4729: out<=1;
   4730: out<=1;
   4731: out<=0;
   4732: out<=0;
   4733: out<=0;
   4734: out<=0;
   4735: out<=0;
   4736: out<=1;
   4737: out<=1;
   4738: out<=0;
   4739: out<=0;
   4740: out<=1;
   4741: out<=0;
   4742: out<=1;
   4743: out<=0;
   4744: out<=1;
   4745: out<=0;
   4746: out<=0;
   4747: out<=1;
   4748: out<=1;
   4749: out<=1;
   4750: out<=1;
   4751: out<=1;
   4752: out<=1;
   4753: out<=1;
   4754: out<=0;
   4755: out<=0;
   4756: out<=1;
   4757: out<=0;
   4758: out<=1;
   4759: out<=0;
   4760: out<=1;
   4761: out<=0;
   4762: out<=0;
   4763: out<=1;
   4764: out<=1;
   4765: out<=1;
   4766: out<=1;
   4767: out<=1;
   4768: out<=0;
   4769: out<=0;
   4770: out<=1;
   4771: out<=1;
   4772: out<=0;
   4773: out<=1;
   4774: out<=0;
   4775: out<=1;
   4776: out<=0;
   4777: out<=1;
   4778: out<=1;
   4779: out<=0;
   4780: out<=0;
   4781: out<=0;
   4782: out<=0;
   4783: out<=0;
   4784: out<=0;
   4785: out<=0;
   4786: out<=1;
   4787: out<=1;
   4788: out<=0;
   4789: out<=1;
   4790: out<=0;
   4791: out<=1;
   4792: out<=0;
   4793: out<=1;
   4794: out<=1;
   4795: out<=0;
   4796: out<=0;
   4797: out<=0;
   4798: out<=0;
   4799: out<=0;
   4800: out<=1;
   4801: out<=1;
   4802: out<=0;
   4803: out<=0;
   4804: out<=1;
   4805: out<=0;
   4806: out<=1;
   4807: out<=0;
   4808: out<=1;
   4809: out<=0;
   4810: out<=0;
   4811: out<=1;
   4812: out<=1;
   4813: out<=1;
   4814: out<=1;
   4815: out<=1;
   4816: out<=0;
   4817: out<=0;
   4818: out<=1;
   4819: out<=1;
   4820: out<=0;
   4821: out<=1;
   4822: out<=0;
   4823: out<=1;
   4824: out<=0;
   4825: out<=1;
   4826: out<=1;
   4827: out<=0;
   4828: out<=0;
   4829: out<=0;
   4830: out<=0;
   4831: out<=0;
   4832: out<=1;
   4833: out<=1;
   4834: out<=0;
   4835: out<=0;
   4836: out<=1;
   4837: out<=0;
   4838: out<=1;
   4839: out<=0;
   4840: out<=1;
   4841: out<=0;
   4842: out<=0;
   4843: out<=1;
   4844: out<=1;
   4845: out<=1;
   4846: out<=1;
   4847: out<=1;
   4848: out<=0;
   4849: out<=0;
   4850: out<=1;
   4851: out<=1;
   4852: out<=0;
   4853: out<=1;
   4854: out<=0;
   4855: out<=1;
   4856: out<=0;
   4857: out<=1;
   4858: out<=1;
   4859: out<=0;
   4860: out<=0;
   4861: out<=0;
   4862: out<=0;
   4863: out<=0;
   4864: out<=0;
   4865: out<=1;
   4866: out<=0;
   4867: out<=1;
   4868: out<=1;
   4869: out<=1;
   4870: out<=0;
   4871: out<=0;
   4872: out<=1;
   4873: out<=1;
   4874: out<=1;
   4875: out<=1;
   4876: out<=0;
   4877: out<=1;
   4878: out<=1;
   4879: out<=0;
   4880: out<=0;
   4881: out<=1;
   4882: out<=0;
   4883: out<=1;
   4884: out<=1;
   4885: out<=1;
   4886: out<=0;
   4887: out<=0;
   4888: out<=1;
   4889: out<=1;
   4890: out<=1;
   4891: out<=1;
   4892: out<=0;
   4893: out<=1;
   4894: out<=1;
   4895: out<=0;
   4896: out<=0;
   4897: out<=1;
   4898: out<=0;
   4899: out<=1;
   4900: out<=1;
   4901: out<=1;
   4902: out<=0;
   4903: out<=0;
   4904: out<=1;
   4905: out<=1;
   4906: out<=1;
   4907: out<=1;
   4908: out<=0;
   4909: out<=1;
   4910: out<=1;
   4911: out<=0;
   4912: out<=0;
   4913: out<=1;
   4914: out<=0;
   4915: out<=1;
   4916: out<=1;
   4917: out<=1;
   4918: out<=0;
   4919: out<=0;
   4920: out<=1;
   4921: out<=1;
   4922: out<=1;
   4923: out<=1;
   4924: out<=0;
   4925: out<=1;
   4926: out<=1;
   4927: out<=0;
   4928: out<=0;
   4929: out<=1;
   4930: out<=0;
   4931: out<=1;
   4932: out<=1;
   4933: out<=1;
   4934: out<=0;
   4935: out<=0;
   4936: out<=1;
   4937: out<=1;
   4938: out<=1;
   4939: out<=1;
   4940: out<=0;
   4941: out<=1;
   4942: out<=1;
   4943: out<=0;
   4944: out<=1;
   4945: out<=0;
   4946: out<=1;
   4947: out<=0;
   4948: out<=0;
   4949: out<=0;
   4950: out<=1;
   4951: out<=1;
   4952: out<=0;
   4953: out<=0;
   4954: out<=0;
   4955: out<=0;
   4956: out<=1;
   4957: out<=0;
   4958: out<=0;
   4959: out<=1;
   4960: out<=1;
   4961: out<=0;
   4962: out<=1;
   4963: out<=0;
   4964: out<=0;
   4965: out<=0;
   4966: out<=1;
   4967: out<=1;
   4968: out<=0;
   4969: out<=0;
   4970: out<=0;
   4971: out<=0;
   4972: out<=1;
   4973: out<=0;
   4974: out<=0;
   4975: out<=1;
   4976: out<=0;
   4977: out<=1;
   4978: out<=0;
   4979: out<=1;
   4980: out<=1;
   4981: out<=1;
   4982: out<=0;
   4983: out<=0;
   4984: out<=1;
   4985: out<=1;
   4986: out<=1;
   4987: out<=1;
   4988: out<=0;
   4989: out<=1;
   4990: out<=1;
   4991: out<=0;
   4992: out<=1;
   4993: out<=0;
   4994: out<=1;
   4995: out<=0;
   4996: out<=0;
   4997: out<=0;
   4998: out<=1;
   4999: out<=1;
   5000: out<=0;
   5001: out<=0;
   5002: out<=0;
   5003: out<=0;
   5004: out<=1;
   5005: out<=0;
   5006: out<=0;
   5007: out<=1;
   5008: out<=0;
   5009: out<=1;
   5010: out<=0;
   5011: out<=1;
   5012: out<=1;
   5013: out<=1;
   5014: out<=0;
   5015: out<=0;
   5016: out<=1;
   5017: out<=1;
   5018: out<=1;
   5019: out<=1;
   5020: out<=0;
   5021: out<=1;
   5022: out<=1;
   5023: out<=0;
   5024: out<=1;
   5025: out<=0;
   5026: out<=1;
   5027: out<=0;
   5028: out<=0;
   5029: out<=0;
   5030: out<=1;
   5031: out<=1;
   5032: out<=0;
   5033: out<=0;
   5034: out<=0;
   5035: out<=0;
   5036: out<=1;
   5037: out<=0;
   5038: out<=0;
   5039: out<=1;
   5040: out<=0;
   5041: out<=1;
   5042: out<=0;
   5043: out<=1;
   5044: out<=1;
   5045: out<=1;
   5046: out<=0;
   5047: out<=0;
   5048: out<=1;
   5049: out<=1;
   5050: out<=1;
   5051: out<=1;
   5052: out<=0;
   5053: out<=1;
   5054: out<=1;
   5055: out<=0;
   5056: out<=1;
   5057: out<=0;
   5058: out<=1;
   5059: out<=0;
   5060: out<=0;
   5061: out<=0;
   5062: out<=1;
   5063: out<=1;
   5064: out<=0;
   5065: out<=0;
   5066: out<=0;
   5067: out<=0;
   5068: out<=1;
   5069: out<=0;
   5070: out<=0;
   5071: out<=1;
   5072: out<=1;
   5073: out<=0;
   5074: out<=1;
   5075: out<=0;
   5076: out<=0;
   5077: out<=0;
   5078: out<=1;
   5079: out<=1;
   5080: out<=0;
   5081: out<=0;
   5082: out<=0;
   5083: out<=0;
   5084: out<=1;
   5085: out<=0;
   5086: out<=0;
   5087: out<=1;
   5088: out<=0;
   5089: out<=1;
   5090: out<=0;
   5091: out<=1;
   5092: out<=1;
   5093: out<=1;
   5094: out<=0;
   5095: out<=0;
   5096: out<=1;
   5097: out<=1;
   5098: out<=1;
   5099: out<=1;
   5100: out<=0;
   5101: out<=1;
   5102: out<=1;
   5103: out<=0;
   5104: out<=0;
   5105: out<=1;
   5106: out<=0;
   5107: out<=1;
   5108: out<=1;
   5109: out<=1;
   5110: out<=0;
   5111: out<=0;
   5112: out<=1;
   5113: out<=1;
   5114: out<=1;
   5115: out<=1;
   5116: out<=0;
   5117: out<=1;
   5118: out<=1;
   5119: out<=0;
   5120: out<=0;
   5121: out<=0;
   5122: out<=0;
   5123: out<=0;
   5124: out<=1;
   5125: out<=0;
   5126: out<=0;
   5127: out<=1;
   5128: out<=0;
   5129: out<=1;
   5130: out<=0;
   5131: out<=1;
   5132: out<=1;
   5133: out<=1;
   5134: out<=0;
   5135: out<=0;
   5136: out<=0;
   5137: out<=0;
   5138: out<=0;
   5139: out<=0;
   5140: out<=1;
   5141: out<=0;
   5142: out<=0;
   5143: out<=1;
   5144: out<=0;
   5145: out<=1;
   5146: out<=0;
   5147: out<=1;
   5148: out<=1;
   5149: out<=1;
   5150: out<=0;
   5151: out<=0;
   5152: out<=1;
   5153: out<=1;
   5154: out<=1;
   5155: out<=1;
   5156: out<=0;
   5157: out<=1;
   5158: out<=1;
   5159: out<=0;
   5160: out<=1;
   5161: out<=0;
   5162: out<=1;
   5163: out<=0;
   5164: out<=0;
   5165: out<=0;
   5166: out<=1;
   5167: out<=1;
   5168: out<=1;
   5169: out<=1;
   5170: out<=1;
   5171: out<=1;
   5172: out<=0;
   5173: out<=1;
   5174: out<=1;
   5175: out<=0;
   5176: out<=1;
   5177: out<=0;
   5178: out<=1;
   5179: out<=0;
   5180: out<=0;
   5181: out<=0;
   5182: out<=1;
   5183: out<=1;
   5184: out<=0;
   5185: out<=0;
   5186: out<=0;
   5187: out<=0;
   5188: out<=1;
   5189: out<=0;
   5190: out<=0;
   5191: out<=1;
   5192: out<=0;
   5193: out<=1;
   5194: out<=0;
   5195: out<=1;
   5196: out<=1;
   5197: out<=1;
   5198: out<=0;
   5199: out<=0;
   5200: out<=1;
   5201: out<=1;
   5202: out<=1;
   5203: out<=1;
   5204: out<=0;
   5205: out<=1;
   5206: out<=1;
   5207: out<=0;
   5208: out<=1;
   5209: out<=0;
   5210: out<=1;
   5211: out<=0;
   5212: out<=0;
   5213: out<=0;
   5214: out<=1;
   5215: out<=1;
   5216: out<=0;
   5217: out<=0;
   5218: out<=0;
   5219: out<=0;
   5220: out<=1;
   5221: out<=0;
   5222: out<=0;
   5223: out<=1;
   5224: out<=0;
   5225: out<=1;
   5226: out<=0;
   5227: out<=1;
   5228: out<=1;
   5229: out<=1;
   5230: out<=0;
   5231: out<=0;
   5232: out<=1;
   5233: out<=1;
   5234: out<=1;
   5235: out<=1;
   5236: out<=0;
   5237: out<=1;
   5238: out<=1;
   5239: out<=0;
   5240: out<=1;
   5241: out<=0;
   5242: out<=1;
   5243: out<=0;
   5244: out<=0;
   5245: out<=0;
   5246: out<=1;
   5247: out<=1;
   5248: out<=1;
   5249: out<=1;
   5250: out<=1;
   5251: out<=1;
   5252: out<=0;
   5253: out<=1;
   5254: out<=1;
   5255: out<=0;
   5256: out<=1;
   5257: out<=0;
   5258: out<=1;
   5259: out<=0;
   5260: out<=0;
   5261: out<=0;
   5262: out<=1;
   5263: out<=1;
   5264: out<=0;
   5265: out<=0;
   5266: out<=0;
   5267: out<=0;
   5268: out<=1;
   5269: out<=0;
   5270: out<=0;
   5271: out<=1;
   5272: out<=0;
   5273: out<=1;
   5274: out<=0;
   5275: out<=1;
   5276: out<=1;
   5277: out<=1;
   5278: out<=0;
   5279: out<=0;
   5280: out<=0;
   5281: out<=0;
   5282: out<=0;
   5283: out<=0;
   5284: out<=1;
   5285: out<=0;
   5286: out<=0;
   5287: out<=1;
   5288: out<=0;
   5289: out<=1;
   5290: out<=0;
   5291: out<=1;
   5292: out<=1;
   5293: out<=1;
   5294: out<=0;
   5295: out<=0;
   5296: out<=1;
   5297: out<=1;
   5298: out<=1;
   5299: out<=1;
   5300: out<=0;
   5301: out<=1;
   5302: out<=1;
   5303: out<=0;
   5304: out<=1;
   5305: out<=0;
   5306: out<=1;
   5307: out<=0;
   5308: out<=0;
   5309: out<=0;
   5310: out<=1;
   5311: out<=1;
   5312: out<=1;
   5313: out<=1;
   5314: out<=1;
   5315: out<=1;
   5316: out<=0;
   5317: out<=1;
   5318: out<=1;
   5319: out<=0;
   5320: out<=1;
   5321: out<=0;
   5322: out<=1;
   5323: out<=0;
   5324: out<=0;
   5325: out<=0;
   5326: out<=1;
   5327: out<=1;
   5328: out<=1;
   5329: out<=1;
   5330: out<=1;
   5331: out<=1;
   5332: out<=0;
   5333: out<=1;
   5334: out<=1;
   5335: out<=0;
   5336: out<=1;
   5337: out<=0;
   5338: out<=1;
   5339: out<=0;
   5340: out<=0;
   5341: out<=0;
   5342: out<=1;
   5343: out<=1;
   5344: out<=1;
   5345: out<=1;
   5346: out<=1;
   5347: out<=1;
   5348: out<=0;
   5349: out<=1;
   5350: out<=1;
   5351: out<=0;
   5352: out<=1;
   5353: out<=0;
   5354: out<=1;
   5355: out<=0;
   5356: out<=0;
   5357: out<=0;
   5358: out<=1;
   5359: out<=1;
   5360: out<=1;
   5361: out<=1;
   5362: out<=1;
   5363: out<=1;
   5364: out<=0;
   5365: out<=1;
   5366: out<=1;
   5367: out<=0;
   5368: out<=1;
   5369: out<=0;
   5370: out<=1;
   5371: out<=0;
   5372: out<=0;
   5373: out<=0;
   5374: out<=1;
   5375: out<=1;
   5376: out<=1;
   5377: out<=0;
   5378: out<=0;
   5379: out<=1;
   5380: out<=1;
   5381: out<=1;
   5382: out<=1;
   5383: out<=1;
   5384: out<=0;
   5385: out<=0;
   5386: out<=1;
   5387: out<=1;
   5388: out<=0;
   5389: out<=1;
   5390: out<=0;
   5391: out<=1;
   5392: out<=0;
   5393: out<=1;
   5394: out<=1;
   5395: out<=0;
   5396: out<=0;
   5397: out<=0;
   5398: out<=0;
   5399: out<=0;
   5400: out<=1;
   5401: out<=1;
   5402: out<=0;
   5403: out<=0;
   5404: out<=1;
   5405: out<=0;
   5406: out<=1;
   5407: out<=0;
   5408: out<=1;
   5409: out<=0;
   5410: out<=0;
   5411: out<=1;
   5412: out<=1;
   5413: out<=1;
   5414: out<=1;
   5415: out<=1;
   5416: out<=0;
   5417: out<=0;
   5418: out<=1;
   5419: out<=1;
   5420: out<=0;
   5421: out<=1;
   5422: out<=0;
   5423: out<=1;
   5424: out<=0;
   5425: out<=1;
   5426: out<=1;
   5427: out<=0;
   5428: out<=0;
   5429: out<=0;
   5430: out<=0;
   5431: out<=0;
   5432: out<=1;
   5433: out<=1;
   5434: out<=0;
   5435: out<=0;
   5436: out<=1;
   5437: out<=0;
   5438: out<=1;
   5439: out<=0;
   5440: out<=1;
   5441: out<=0;
   5442: out<=0;
   5443: out<=1;
   5444: out<=1;
   5445: out<=1;
   5446: out<=1;
   5447: out<=1;
   5448: out<=0;
   5449: out<=0;
   5450: out<=1;
   5451: out<=1;
   5452: out<=0;
   5453: out<=1;
   5454: out<=0;
   5455: out<=1;
   5456: out<=1;
   5457: out<=0;
   5458: out<=0;
   5459: out<=1;
   5460: out<=1;
   5461: out<=1;
   5462: out<=1;
   5463: out<=1;
   5464: out<=0;
   5465: out<=0;
   5466: out<=1;
   5467: out<=1;
   5468: out<=0;
   5469: out<=1;
   5470: out<=0;
   5471: out<=1;
   5472: out<=0;
   5473: out<=1;
   5474: out<=1;
   5475: out<=0;
   5476: out<=0;
   5477: out<=0;
   5478: out<=0;
   5479: out<=0;
   5480: out<=1;
   5481: out<=1;
   5482: out<=0;
   5483: out<=0;
   5484: out<=1;
   5485: out<=0;
   5486: out<=1;
   5487: out<=0;
   5488: out<=0;
   5489: out<=1;
   5490: out<=1;
   5491: out<=0;
   5492: out<=0;
   5493: out<=0;
   5494: out<=0;
   5495: out<=0;
   5496: out<=1;
   5497: out<=1;
   5498: out<=0;
   5499: out<=0;
   5500: out<=1;
   5501: out<=0;
   5502: out<=1;
   5503: out<=0;
   5504: out<=0;
   5505: out<=1;
   5506: out<=1;
   5507: out<=0;
   5508: out<=0;
   5509: out<=0;
   5510: out<=0;
   5511: out<=0;
   5512: out<=1;
   5513: out<=1;
   5514: out<=0;
   5515: out<=0;
   5516: out<=1;
   5517: out<=0;
   5518: out<=1;
   5519: out<=0;
   5520: out<=0;
   5521: out<=1;
   5522: out<=1;
   5523: out<=0;
   5524: out<=0;
   5525: out<=0;
   5526: out<=0;
   5527: out<=0;
   5528: out<=1;
   5529: out<=1;
   5530: out<=0;
   5531: out<=0;
   5532: out<=1;
   5533: out<=0;
   5534: out<=1;
   5535: out<=0;
   5536: out<=0;
   5537: out<=1;
   5538: out<=1;
   5539: out<=0;
   5540: out<=0;
   5541: out<=0;
   5542: out<=0;
   5543: out<=0;
   5544: out<=1;
   5545: out<=1;
   5546: out<=0;
   5547: out<=0;
   5548: out<=1;
   5549: out<=0;
   5550: out<=1;
   5551: out<=0;
   5552: out<=0;
   5553: out<=1;
   5554: out<=1;
   5555: out<=0;
   5556: out<=0;
   5557: out<=0;
   5558: out<=0;
   5559: out<=0;
   5560: out<=1;
   5561: out<=1;
   5562: out<=0;
   5563: out<=0;
   5564: out<=1;
   5565: out<=0;
   5566: out<=1;
   5567: out<=0;
   5568: out<=0;
   5569: out<=1;
   5570: out<=1;
   5571: out<=0;
   5572: out<=0;
   5573: out<=0;
   5574: out<=0;
   5575: out<=0;
   5576: out<=1;
   5577: out<=1;
   5578: out<=0;
   5579: out<=0;
   5580: out<=1;
   5581: out<=0;
   5582: out<=1;
   5583: out<=0;
   5584: out<=1;
   5585: out<=0;
   5586: out<=0;
   5587: out<=1;
   5588: out<=1;
   5589: out<=1;
   5590: out<=1;
   5591: out<=1;
   5592: out<=0;
   5593: out<=0;
   5594: out<=1;
   5595: out<=1;
   5596: out<=0;
   5597: out<=1;
   5598: out<=0;
   5599: out<=1;
   5600: out<=1;
   5601: out<=0;
   5602: out<=0;
   5603: out<=1;
   5604: out<=1;
   5605: out<=1;
   5606: out<=1;
   5607: out<=1;
   5608: out<=0;
   5609: out<=0;
   5610: out<=1;
   5611: out<=1;
   5612: out<=0;
   5613: out<=1;
   5614: out<=0;
   5615: out<=1;
   5616: out<=0;
   5617: out<=1;
   5618: out<=1;
   5619: out<=0;
   5620: out<=0;
   5621: out<=0;
   5622: out<=0;
   5623: out<=0;
   5624: out<=1;
   5625: out<=1;
   5626: out<=0;
   5627: out<=0;
   5628: out<=1;
   5629: out<=0;
   5630: out<=1;
   5631: out<=0;
   5632: out<=1;
   5633: out<=0;
   5634: out<=1;
   5635: out<=0;
   5636: out<=1;
   5637: out<=1;
   5638: out<=0;
   5639: out<=0;
   5640: out<=1;
   5641: out<=1;
   5642: out<=1;
   5643: out<=1;
   5644: out<=1;
   5645: out<=0;
   5646: out<=0;
   5647: out<=1;
   5648: out<=0;
   5649: out<=1;
   5650: out<=0;
   5651: out<=1;
   5652: out<=0;
   5653: out<=0;
   5654: out<=1;
   5655: out<=1;
   5656: out<=0;
   5657: out<=0;
   5658: out<=0;
   5659: out<=0;
   5660: out<=0;
   5661: out<=1;
   5662: out<=1;
   5663: out<=0;
   5664: out<=0;
   5665: out<=1;
   5666: out<=0;
   5667: out<=1;
   5668: out<=0;
   5669: out<=0;
   5670: out<=1;
   5671: out<=1;
   5672: out<=0;
   5673: out<=0;
   5674: out<=0;
   5675: out<=0;
   5676: out<=0;
   5677: out<=1;
   5678: out<=1;
   5679: out<=0;
   5680: out<=1;
   5681: out<=0;
   5682: out<=1;
   5683: out<=0;
   5684: out<=1;
   5685: out<=1;
   5686: out<=0;
   5687: out<=0;
   5688: out<=1;
   5689: out<=1;
   5690: out<=1;
   5691: out<=1;
   5692: out<=1;
   5693: out<=0;
   5694: out<=0;
   5695: out<=1;
   5696: out<=1;
   5697: out<=0;
   5698: out<=1;
   5699: out<=0;
   5700: out<=1;
   5701: out<=1;
   5702: out<=0;
   5703: out<=0;
   5704: out<=1;
   5705: out<=1;
   5706: out<=1;
   5707: out<=1;
   5708: out<=1;
   5709: out<=0;
   5710: out<=0;
   5711: out<=1;
   5712: out<=1;
   5713: out<=0;
   5714: out<=1;
   5715: out<=0;
   5716: out<=1;
   5717: out<=1;
   5718: out<=0;
   5719: out<=0;
   5720: out<=1;
   5721: out<=1;
   5722: out<=1;
   5723: out<=1;
   5724: out<=1;
   5725: out<=0;
   5726: out<=0;
   5727: out<=1;
   5728: out<=1;
   5729: out<=0;
   5730: out<=1;
   5731: out<=0;
   5732: out<=1;
   5733: out<=1;
   5734: out<=0;
   5735: out<=0;
   5736: out<=1;
   5737: out<=1;
   5738: out<=1;
   5739: out<=1;
   5740: out<=1;
   5741: out<=0;
   5742: out<=0;
   5743: out<=1;
   5744: out<=1;
   5745: out<=0;
   5746: out<=1;
   5747: out<=0;
   5748: out<=1;
   5749: out<=1;
   5750: out<=0;
   5751: out<=0;
   5752: out<=1;
   5753: out<=1;
   5754: out<=1;
   5755: out<=1;
   5756: out<=1;
   5757: out<=0;
   5758: out<=0;
   5759: out<=1;
   5760: out<=0;
   5761: out<=1;
   5762: out<=0;
   5763: out<=1;
   5764: out<=0;
   5765: out<=0;
   5766: out<=1;
   5767: out<=1;
   5768: out<=0;
   5769: out<=0;
   5770: out<=0;
   5771: out<=0;
   5772: out<=0;
   5773: out<=1;
   5774: out<=1;
   5775: out<=0;
   5776: out<=0;
   5777: out<=1;
   5778: out<=0;
   5779: out<=1;
   5780: out<=0;
   5781: out<=0;
   5782: out<=1;
   5783: out<=1;
   5784: out<=0;
   5785: out<=0;
   5786: out<=0;
   5787: out<=0;
   5788: out<=0;
   5789: out<=1;
   5790: out<=1;
   5791: out<=0;
   5792: out<=1;
   5793: out<=0;
   5794: out<=1;
   5795: out<=0;
   5796: out<=1;
   5797: out<=1;
   5798: out<=0;
   5799: out<=0;
   5800: out<=1;
   5801: out<=1;
   5802: out<=1;
   5803: out<=1;
   5804: out<=1;
   5805: out<=0;
   5806: out<=0;
   5807: out<=1;
   5808: out<=1;
   5809: out<=0;
   5810: out<=1;
   5811: out<=0;
   5812: out<=1;
   5813: out<=1;
   5814: out<=0;
   5815: out<=0;
   5816: out<=1;
   5817: out<=1;
   5818: out<=1;
   5819: out<=1;
   5820: out<=1;
   5821: out<=0;
   5822: out<=0;
   5823: out<=1;
   5824: out<=0;
   5825: out<=1;
   5826: out<=0;
   5827: out<=1;
   5828: out<=0;
   5829: out<=0;
   5830: out<=1;
   5831: out<=1;
   5832: out<=0;
   5833: out<=0;
   5834: out<=0;
   5835: out<=0;
   5836: out<=0;
   5837: out<=1;
   5838: out<=1;
   5839: out<=0;
   5840: out<=1;
   5841: out<=0;
   5842: out<=1;
   5843: out<=0;
   5844: out<=1;
   5845: out<=1;
   5846: out<=0;
   5847: out<=0;
   5848: out<=1;
   5849: out<=1;
   5850: out<=1;
   5851: out<=1;
   5852: out<=1;
   5853: out<=0;
   5854: out<=0;
   5855: out<=1;
   5856: out<=0;
   5857: out<=1;
   5858: out<=0;
   5859: out<=1;
   5860: out<=0;
   5861: out<=0;
   5862: out<=1;
   5863: out<=1;
   5864: out<=0;
   5865: out<=0;
   5866: out<=0;
   5867: out<=0;
   5868: out<=0;
   5869: out<=1;
   5870: out<=1;
   5871: out<=0;
   5872: out<=1;
   5873: out<=0;
   5874: out<=1;
   5875: out<=0;
   5876: out<=1;
   5877: out<=1;
   5878: out<=0;
   5879: out<=0;
   5880: out<=1;
   5881: out<=1;
   5882: out<=1;
   5883: out<=1;
   5884: out<=1;
   5885: out<=0;
   5886: out<=0;
   5887: out<=1;
   5888: out<=0;
   5889: out<=0;
   5890: out<=1;
   5891: out<=1;
   5892: out<=1;
   5893: out<=0;
   5894: out<=1;
   5895: out<=0;
   5896: out<=1;
   5897: out<=0;
   5898: out<=0;
   5899: out<=1;
   5900: out<=0;
   5901: out<=0;
   5902: out<=0;
   5903: out<=0;
   5904: out<=0;
   5905: out<=0;
   5906: out<=1;
   5907: out<=1;
   5908: out<=1;
   5909: out<=0;
   5910: out<=1;
   5911: out<=0;
   5912: out<=1;
   5913: out<=0;
   5914: out<=0;
   5915: out<=1;
   5916: out<=0;
   5917: out<=0;
   5918: out<=0;
   5919: out<=0;
   5920: out<=0;
   5921: out<=0;
   5922: out<=1;
   5923: out<=1;
   5924: out<=1;
   5925: out<=0;
   5926: out<=1;
   5927: out<=0;
   5928: out<=1;
   5929: out<=0;
   5930: out<=0;
   5931: out<=1;
   5932: out<=0;
   5933: out<=0;
   5934: out<=0;
   5935: out<=0;
   5936: out<=0;
   5937: out<=0;
   5938: out<=1;
   5939: out<=1;
   5940: out<=1;
   5941: out<=0;
   5942: out<=1;
   5943: out<=0;
   5944: out<=1;
   5945: out<=0;
   5946: out<=0;
   5947: out<=1;
   5948: out<=0;
   5949: out<=0;
   5950: out<=0;
   5951: out<=0;
   5952: out<=0;
   5953: out<=0;
   5954: out<=1;
   5955: out<=1;
   5956: out<=1;
   5957: out<=0;
   5958: out<=1;
   5959: out<=0;
   5960: out<=1;
   5961: out<=0;
   5962: out<=0;
   5963: out<=1;
   5964: out<=0;
   5965: out<=0;
   5966: out<=0;
   5967: out<=0;
   5968: out<=1;
   5969: out<=1;
   5970: out<=0;
   5971: out<=0;
   5972: out<=0;
   5973: out<=1;
   5974: out<=0;
   5975: out<=1;
   5976: out<=0;
   5977: out<=1;
   5978: out<=1;
   5979: out<=0;
   5980: out<=1;
   5981: out<=1;
   5982: out<=1;
   5983: out<=1;
   5984: out<=1;
   5985: out<=1;
   5986: out<=0;
   5987: out<=0;
   5988: out<=0;
   5989: out<=1;
   5990: out<=0;
   5991: out<=1;
   5992: out<=0;
   5993: out<=1;
   5994: out<=1;
   5995: out<=0;
   5996: out<=1;
   5997: out<=1;
   5998: out<=1;
   5999: out<=1;
   6000: out<=0;
   6001: out<=0;
   6002: out<=1;
   6003: out<=1;
   6004: out<=1;
   6005: out<=0;
   6006: out<=1;
   6007: out<=0;
   6008: out<=1;
   6009: out<=0;
   6010: out<=0;
   6011: out<=1;
   6012: out<=0;
   6013: out<=0;
   6014: out<=0;
   6015: out<=0;
   6016: out<=1;
   6017: out<=1;
   6018: out<=0;
   6019: out<=0;
   6020: out<=0;
   6021: out<=1;
   6022: out<=0;
   6023: out<=1;
   6024: out<=0;
   6025: out<=1;
   6026: out<=1;
   6027: out<=0;
   6028: out<=1;
   6029: out<=1;
   6030: out<=1;
   6031: out<=1;
   6032: out<=0;
   6033: out<=0;
   6034: out<=1;
   6035: out<=1;
   6036: out<=1;
   6037: out<=0;
   6038: out<=1;
   6039: out<=0;
   6040: out<=1;
   6041: out<=0;
   6042: out<=0;
   6043: out<=1;
   6044: out<=0;
   6045: out<=0;
   6046: out<=0;
   6047: out<=0;
   6048: out<=1;
   6049: out<=1;
   6050: out<=0;
   6051: out<=0;
   6052: out<=0;
   6053: out<=1;
   6054: out<=0;
   6055: out<=1;
   6056: out<=0;
   6057: out<=1;
   6058: out<=1;
   6059: out<=0;
   6060: out<=1;
   6061: out<=1;
   6062: out<=1;
   6063: out<=1;
   6064: out<=0;
   6065: out<=0;
   6066: out<=1;
   6067: out<=1;
   6068: out<=1;
   6069: out<=0;
   6070: out<=1;
   6071: out<=0;
   6072: out<=1;
   6073: out<=0;
   6074: out<=0;
   6075: out<=1;
   6076: out<=0;
   6077: out<=0;
   6078: out<=0;
   6079: out<=0;
   6080: out<=1;
   6081: out<=1;
   6082: out<=0;
   6083: out<=0;
   6084: out<=0;
   6085: out<=1;
   6086: out<=0;
   6087: out<=1;
   6088: out<=0;
   6089: out<=1;
   6090: out<=1;
   6091: out<=0;
   6092: out<=1;
   6093: out<=1;
   6094: out<=1;
   6095: out<=1;
   6096: out<=1;
   6097: out<=1;
   6098: out<=0;
   6099: out<=0;
   6100: out<=0;
   6101: out<=1;
   6102: out<=0;
   6103: out<=1;
   6104: out<=0;
   6105: out<=1;
   6106: out<=1;
   6107: out<=0;
   6108: out<=1;
   6109: out<=1;
   6110: out<=1;
   6111: out<=1;
   6112: out<=0;
   6113: out<=0;
   6114: out<=1;
   6115: out<=1;
   6116: out<=1;
   6117: out<=0;
   6118: out<=1;
   6119: out<=0;
   6120: out<=1;
   6121: out<=0;
   6122: out<=0;
   6123: out<=1;
   6124: out<=0;
   6125: out<=0;
   6126: out<=0;
   6127: out<=0;
   6128: out<=0;
   6129: out<=0;
   6130: out<=1;
   6131: out<=1;
   6132: out<=1;
   6133: out<=0;
   6134: out<=1;
   6135: out<=0;
   6136: out<=1;
   6137: out<=0;
   6138: out<=0;
   6139: out<=1;
   6140: out<=0;
   6141: out<=0;
   6142: out<=0;
   6143: out<=0;
   6144: out<=0;
   6145: out<=0;
   6146: out<=1;
   6147: out<=1;
   6148: out<=1;
   6149: out<=0;
   6150: out<=1;
   6151: out<=0;
   6152: out<=0;
   6153: out<=1;
   6154: out<=1;
   6155: out<=0;
   6156: out<=1;
   6157: out<=1;
   6158: out<=1;
   6159: out<=1;
   6160: out<=0;
   6161: out<=0;
   6162: out<=1;
   6163: out<=1;
   6164: out<=1;
   6165: out<=0;
   6166: out<=1;
   6167: out<=0;
   6168: out<=0;
   6169: out<=1;
   6170: out<=1;
   6171: out<=0;
   6172: out<=1;
   6173: out<=1;
   6174: out<=1;
   6175: out<=1;
   6176: out<=1;
   6177: out<=1;
   6178: out<=0;
   6179: out<=0;
   6180: out<=0;
   6181: out<=1;
   6182: out<=0;
   6183: out<=1;
   6184: out<=1;
   6185: out<=0;
   6186: out<=0;
   6187: out<=1;
   6188: out<=0;
   6189: out<=0;
   6190: out<=0;
   6191: out<=0;
   6192: out<=1;
   6193: out<=1;
   6194: out<=0;
   6195: out<=0;
   6196: out<=0;
   6197: out<=1;
   6198: out<=0;
   6199: out<=1;
   6200: out<=1;
   6201: out<=0;
   6202: out<=0;
   6203: out<=1;
   6204: out<=0;
   6205: out<=0;
   6206: out<=0;
   6207: out<=0;
   6208: out<=0;
   6209: out<=0;
   6210: out<=1;
   6211: out<=1;
   6212: out<=1;
   6213: out<=0;
   6214: out<=1;
   6215: out<=0;
   6216: out<=0;
   6217: out<=1;
   6218: out<=1;
   6219: out<=0;
   6220: out<=1;
   6221: out<=1;
   6222: out<=1;
   6223: out<=1;
   6224: out<=1;
   6225: out<=1;
   6226: out<=0;
   6227: out<=0;
   6228: out<=0;
   6229: out<=1;
   6230: out<=0;
   6231: out<=1;
   6232: out<=1;
   6233: out<=0;
   6234: out<=0;
   6235: out<=1;
   6236: out<=0;
   6237: out<=0;
   6238: out<=0;
   6239: out<=0;
   6240: out<=0;
   6241: out<=0;
   6242: out<=1;
   6243: out<=1;
   6244: out<=1;
   6245: out<=0;
   6246: out<=1;
   6247: out<=0;
   6248: out<=0;
   6249: out<=1;
   6250: out<=1;
   6251: out<=0;
   6252: out<=1;
   6253: out<=1;
   6254: out<=1;
   6255: out<=1;
   6256: out<=1;
   6257: out<=1;
   6258: out<=0;
   6259: out<=0;
   6260: out<=0;
   6261: out<=1;
   6262: out<=0;
   6263: out<=1;
   6264: out<=1;
   6265: out<=0;
   6266: out<=0;
   6267: out<=1;
   6268: out<=0;
   6269: out<=0;
   6270: out<=0;
   6271: out<=0;
   6272: out<=1;
   6273: out<=1;
   6274: out<=0;
   6275: out<=0;
   6276: out<=0;
   6277: out<=1;
   6278: out<=0;
   6279: out<=1;
   6280: out<=1;
   6281: out<=0;
   6282: out<=0;
   6283: out<=1;
   6284: out<=0;
   6285: out<=0;
   6286: out<=0;
   6287: out<=0;
   6288: out<=0;
   6289: out<=0;
   6290: out<=1;
   6291: out<=1;
   6292: out<=1;
   6293: out<=0;
   6294: out<=1;
   6295: out<=0;
   6296: out<=0;
   6297: out<=1;
   6298: out<=1;
   6299: out<=0;
   6300: out<=1;
   6301: out<=1;
   6302: out<=1;
   6303: out<=1;
   6304: out<=0;
   6305: out<=0;
   6306: out<=1;
   6307: out<=1;
   6308: out<=1;
   6309: out<=0;
   6310: out<=1;
   6311: out<=0;
   6312: out<=0;
   6313: out<=1;
   6314: out<=1;
   6315: out<=0;
   6316: out<=1;
   6317: out<=1;
   6318: out<=1;
   6319: out<=1;
   6320: out<=1;
   6321: out<=1;
   6322: out<=0;
   6323: out<=0;
   6324: out<=0;
   6325: out<=1;
   6326: out<=0;
   6327: out<=1;
   6328: out<=1;
   6329: out<=0;
   6330: out<=0;
   6331: out<=1;
   6332: out<=0;
   6333: out<=0;
   6334: out<=0;
   6335: out<=0;
   6336: out<=1;
   6337: out<=1;
   6338: out<=0;
   6339: out<=0;
   6340: out<=0;
   6341: out<=1;
   6342: out<=0;
   6343: out<=1;
   6344: out<=1;
   6345: out<=0;
   6346: out<=0;
   6347: out<=1;
   6348: out<=0;
   6349: out<=0;
   6350: out<=0;
   6351: out<=0;
   6352: out<=1;
   6353: out<=1;
   6354: out<=0;
   6355: out<=0;
   6356: out<=0;
   6357: out<=1;
   6358: out<=0;
   6359: out<=1;
   6360: out<=1;
   6361: out<=0;
   6362: out<=0;
   6363: out<=1;
   6364: out<=0;
   6365: out<=0;
   6366: out<=0;
   6367: out<=0;
   6368: out<=1;
   6369: out<=1;
   6370: out<=0;
   6371: out<=0;
   6372: out<=0;
   6373: out<=1;
   6374: out<=0;
   6375: out<=1;
   6376: out<=1;
   6377: out<=0;
   6378: out<=0;
   6379: out<=1;
   6380: out<=0;
   6381: out<=0;
   6382: out<=0;
   6383: out<=0;
   6384: out<=1;
   6385: out<=1;
   6386: out<=0;
   6387: out<=0;
   6388: out<=0;
   6389: out<=1;
   6390: out<=0;
   6391: out<=1;
   6392: out<=1;
   6393: out<=0;
   6394: out<=0;
   6395: out<=1;
   6396: out<=0;
   6397: out<=0;
   6398: out<=0;
   6399: out<=0;
   6400: out<=1;
   6401: out<=0;
   6402: out<=1;
   6403: out<=0;
   6404: out<=1;
   6405: out<=1;
   6406: out<=0;
   6407: out<=0;
   6408: out<=0;
   6409: out<=0;
   6410: out<=0;
   6411: out<=0;
   6412: out<=0;
   6413: out<=1;
   6414: out<=1;
   6415: out<=0;
   6416: out<=0;
   6417: out<=1;
   6418: out<=0;
   6419: out<=1;
   6420: out<=0;
   6421: out<=0;
   6422: out<=1;
   6423: out<=1;
   6424: out<=1;
   6425: out<=1;
   6426: out<=1;
   6427: out<=1;
   6428: out<=1;
   6429: out<=0;
   6430: out<=0;
   6431: out<=1;
   6432: out<=1;
   6433: out<=0;
   6434: out<=1;
   6435: out<=0;
   6436: out<=1;
   6437: out<=1;
   6438: out<=0;
   6439: out<=0;
   6440: out<=0;
   6441: out<=0;
   6442: out<=0;
   6443: out<=0;
   6444: out<=0;
   6445: out<=1;
   6446: out<=1;
   6447: out<=0;
   6448: out<=0;
   6449: out<=1;
   6450: out<=0;
   6451: out<=1;
   6452: out<=0;
   6453: out<=0;
   6454: out<=1;
   6455: out<=1;
   6456: out<=1;
   6457: out<=1;
   6458: out<=1;
   6459: out<=1;
   6460: out<=1;
   6461: out<=0;
   6462: out<=0;
   6463: out<=1;
   6464: out<=1;
   6465: out<=0;
   6466: out<=1;
   6467: out<=0;
   6468: out<=1;
   6469: out<=1;
   6470: out<=0;
   6471: out<=0;
   6472: out<=0;
   6473: out<=0;
   6474: out<=0;
   6475: out<=0;
   6476: out<=0;
   6477: out<=1;
   6478: out<=1;
   6479: out<=0;
   6480: out<=1;
   6481: out<=0;
   6482: out<=1;
   6483: out<=0;
   6484: out<=1;
   6485: out<=1;
   6486: out<=0;
   6487: out<=0;
   6488: out<=0;
   6489: out<=0;
   6490: out<=0;
   6491: out<=0;
   6492: out<=0;
   6493: out<=1;
   6494: out<=1;
   6495: out<=0;
   6496: out<=0;
   6497: out<=1;
   6498: out<=0;
   6499: out<=1;
   6500: out<=0;
   6501: out<=0;
   6502: out<=1;
   6503: out<=1;
   6504: out<=1;
   6505: out<=1;
   6506: out<=1;
   6507: out<=1;
   6508: out<=1;
   6509: out<=0;
   6510: out<=0;
   6511: out<=1;
   6512: out<=0;
   6513: out<=1;
   6514: out<=0;
   6515: out<=1;
   6516: out<=0;
   6517: out<=0;
   6518: out<=1;
   6519: out<=1;
   6520: out<=1;
   6521: out<=1;
   6522: out<=1;
   6523: out<=1;
   6524: out<=1;
   6525: out<=0;
   6526: out<=0;
   6527: out<=1;
   6528: out<=0;
   6529: out<=1;
   6530: out<=0;
   6531: out<=1;
   6532: out<=0;
   6533: out<=0;
   6534: out<=1;
   6535: out<=1;
   6536: out<=1;
   6537: out<=1;
   6538: out<=1;
   6539: out<=1;
   6540: out<=1;
   6541: out<=0;
   6542: out<=0;
   6543: out<=1;
   6544: out<=0;
   6545: out<=1;
   6546: out<=0;
   6547: out<=1;
   6548: out<=0;
   6549: out<=0;
   6550: out<=1;
   6551: out<=1;
   6552: out<=1;
   6553: out<=1;
   6554: out<=1;
   6555: out<=1;
   6556: out<=1;
   6557: out<=0;
   6558: out<=0;
   6559: out<=1;
   6560: out<=0;
   6561: out<=1;
   6562: out<=0;
   6563: out<=1;
   6564: out<=0;
   6565: out<=0;
   6566: out<=1;
   6567: out<=1;
   6568: out<=1;
   6569: out<=1;
   6570: out<=1;
   6571: out<=1;
   6572: out<=1;
   6573: out<=0;
   6574: out<=0;
   6575: out<=1;
   6576: out<=0;
   6577: out<=1;
   6578: out<=0;
   6579: out<=1;
   6580: out<=0;
   6581: out<=0;
   6582: out<=1;
   6583: out<=1;
   6584: out<=1;
   6585: out<=1;
   6586: out<=1;
   6587: out<=1;
   6588: out<=1;
   6589: out<=0;
   6590: out<=0;
   6591: out<=1;
   6592: out<=0;
   6593: out<=1;
   6594: out<=0;
   6595: out<=1;
   6596: out<=0;
   6597: out<=0;
   6598: out<=1;
   6599: out<=1;
   6600: out<=1;
   6601: out<=1;
   6602: out<=1;
   6603: out<=1;
   6604: out<=1;
   6605: out<=0;
   6606: out<=0;
   6607: out<=1;
   6608: out<=1;
   6609: out<=0;
   6610: out<=1;
   6611: out<=0;
   6612: out<=1;
   6613: out<=1;
   6614: out<=0;
   6615: out<=0;
   6616: out<=0;
   6617: out<=0;
   6618: out<=0;
   6619: out<=0;
   6620: out<=0;
   6621: out<=1;
   6622: out<=1;
   6623: out<=0;
   6624: out<=1;
   6625: out<=0;
   6626: out<=1;
   6627: out<=0;
   6628: out<=1;
   6629: out<=1;
   6630: out<=0;
   6631: out<=0;
   6632: out<=0;
   6633: out<=0;
   6634: out<=0;
   6635: out<=0;
   6636: out<=0;
   6637: out<=1;
   6638: out<=1;
   6639: out<=0;
   6640: out<=0;
   6641: out<=1;
   6642: out<=0;
   6643: out<=1;
   6644: out<=0;
   6645: out<=0;
   6646: out<=1;
   6647: out<=1;
   6648: out<=1;
   6649: out<=1;
   6650: out<=1;
   6651: out<=1;
   6652: out<=1;
   6653: out<=0;
   6654: out<=0;
   6655: out<=1;
   6656: out<=0;
   6657: out<=1;
   6658: out<=1;
   6659: out<=0;
   6660: out<=0;
   6661: out<=0;
   6662: out<=0;
   6663: out<=0;
   6664: out<=0;
   6665: out<=0;
   6666: out<=1;
   6667: out<=1;
   6668: out<=0;
   6669: out<=1;
   6670: out<=0;
   6671: out<=1;
   6672: out<=1;
   6673: out<=0;
   6674: out<=0;
   6675: out<=1;
   6676: out<=1;
   6677: out<=1;
   6678: out<=1;
   6679: out<=1;
   6680: out<=1;
   6681: out<=1;
   6682: out<=0;
   6683: out<=0;
   6684: out<=1;
   6685: out<=0;
   6686: out<=1;
   6687: out<=0;
   6688: out<=1;
   6689: out<=0;
   6690: out<=0;
   6691: out<=1;
   6692: out<=1;
   6693: out<=1;
   6694: out<=1;
   6695: out<=1;
   6696: out<=1;
   6697: out<=1;
   6698: out<=0;
   6699: out<=0;
   6700: out<=1;
   6701: out<=0;
   6702: out<=1;
   6703: out<=0;
   6704: out<=0;
   6705: out<=1;
   6706: out<=1;
   6707: out<=0;
   6708: out<=0;
   6709: out<=0;
   6710: out<=0;
   6711: out<=0;
   6712: out<=0;
   6713: out<=0;
   6714: out<=1;
   6715: out<=1;
   6716: out<=0;
   6717: out<=1;
   6718: out<=0;
   6719: out<=1;
   6720: out<=0;
   6721: out<=1;
   6722: out<=1;
   6723: out<=0;
   6724: out<=0;
   6725: out<=0;
   6726: out<=0;
   6727: out<=0;
   6728: out<=0;
   6729: out<=0;
   6730: out<=1;
   6731: out<=1;
   6732: out<=0;
   6733: out<=1;
   6734: out<=0;
   6735: out<=1;
   6736: out<=0;
   6737: out<=1;
   6738: out<=1;
   6739: out<=0;
   6740: out<=0;
   6741: out<=0;
   6742: out<=0;
   6743: out<=0;
   6744: out<=0;
   6745: out<=0;
   6746: out<=1;
   6747: out<=1;
   6748: out<=0;
   6749: out<=1;
   6750: out<=0;
   6751: out<=1;
   6752: out<=0;
   6753: out<=1;
   6754: out<=1;
   6755: out<=0;
   6756: out<=0;
   6757: out<=0;
   6758: out<=0;
   6759: out<=0;
   6760: out<=0;
   6761: out<=0;
   6762: out<=1;
   6763: out<=1;
   6764: out<=0;
   6765: out<=1;
   6766: out<=0;
   6767: out<=1;
   6768: out<=0;
   6769: out<=1;
   6770: out<=1;
   6771: out<=0;
   6772: out<=0;
   6773: out<=0;
   6774: out<=0;
   6775: out<=0;
   6776: out<=0;
   6777: out<=0;
   6778: out<=1;
   6779: out<=1;
   6780: out<=0;
   6781: out<=1;
   6782: out<=0;
   6783: out<=1;
   6784: out<=1;
   6785: out<=0;
   6786: out<=0;
   6787: out<=1;
   6788: out<=1;
   6789: out<=1;
   6790: out<=1;
   6791: out<=1;
   6792: out<=1;
   6793: out<=1;
   6794: out<=0;
   6795: out<=0;
   6796: out<=1;
   6797: out<=0;
   6798: out<=1;
   6799: out<=0;
   6800: out<=1;
   6801: out<=0;
   6802: out<=0;
   6803: out<=1;
   6804: out<=1;
   6805: out<=1;
   6806: out<=1;
   6807: out<=1;
   6808: out<=1;
   6809: out<=1;
   6810: out<=0;
   6811: out<=0;
   6812: out<=1;
   6813: out<=0;
   6814: out<=1;
   6815: out<=0;
   6816: out<=0;
   6817: out<=1;
   6818: out<=1;
   6819: out<=0;
   6820: out<=0;
   6821: out<=0;
   6822: out<=0;
   6823: out<=0;
   6824: out<=0;
   6825: out<=0;
   6826: out<=1;
   6827: out<=1;
   6828: out<=0;
   6829: out<=1;
   6830: out<=0;
   6831: out<=1;
   6832: out<=0;
   6833: out<=1;
   6834: out<=1;
   6835: out<=0;
   6836: out<=0;
   6837: out<=0;
   6838: out<=0;
   6839: out<=0;
   6840: out<=0;
   6841: out<=0;
   6842: out<=1;
   6843: out<=1;
   6844: out<=0;
   6845: out<=1;
   6846: out<=0;
   6847: out<=1;
   6848: out<=1;
   6849: out<=0;
   6850: out<=0;
   6851: out<=1;
   6852: out<=1;
   6853: out<=1;
   6854: out<=1;
   6855: out<=1;
   6856: out<=1;
   6857: out<=1;
   6858: out<=0;
   6859: out<=0;
   6860: out<=1;
   6861: out<=0;
   6862: out<=1;
   6863: out<=0;
   6864: out<=0;
   6865: out<=1;
   6866: out<=1;
   6867: out<=0;
   6868: out<=0;
   6869: out<=0;
   6870: out<=0;
   6871: out<=0;
   6872: out<=0;
   6873: out<=0;
   6874: out<=1;
   6875: out<=1;
   6876: out<=0;
   6877: out<=1;
   6878: out<=0;
   6879: out<=1;
   6880: out<=1;
   6881: out<=0;
   6882: out<=0;
   6883: out<=1;
   6884: out<=1;
   6885: out<=1;
   6886: out<=1;
   6887: out<=1;
   6888: out<=1;
   6889: out<=1;
   6890: out<=0;
   6891: out<=0;
   6892: out<=1;
   6893: out<=0;
   6894: out<=1;
   6895: out<=0;
   6896: out<=0;
   6897: out<=1;
   6898: out<=1;
   6899: out<=0;
   6900: out<=0;
   6901: out<=0;
   6902: out<=0;
   6903: out<=0;
   6904: out<=0;
   6905: out<=0;
   6906: out<=1;
   6907: out<=1;
   6908: out<=0;
   6909: out<=1;
   6910: out<=0;
   6911: out<=1;
   6912: out<=1;
   6913: out<=1;
   6914: out<=1;
   6915: out<=1;
   6916: out<=0;
   6917: out<=1;
   6918: out<=1;
   6919: out<=0;
   6920: out<=0;
   6921: out<=1;
   6922: out<=0;
   6923: out<=1;
   6924: out<=1;
   6925: out<=1;
   6926: out<=0;
   6927: out<=0;
   6928: out<=1;
   6929: out<=1;
   6930: out<=1;
   6931: out<=1;
   6932: out<=0;
   6933: out<=1;
   6934: out<=1;
   6935: out<=0;
   6936: out<=0;
   6937: out<=1;
   6938: out<=0;
   6939: out<=1;
   6940: out<=1;
   6941: out<=1;
   6942: out<=0;
   6943: out<=0;
   6944: out<=1;
   6945: out<=1;
   6946: out<=1;
   6947: out<=1;
   6948: out<=0;
   6949: out<=1;
   6950: out<=1;
   6951: out<=0;
   6952: out<=0;
   6953: out<=1;
   6954: out<=0;
   6955: out<=1;
   6956: out<=1;
   6957: out<=1;
   6958: out<=0;
   6959: out<=0;
   6960: out<=1;
   6961: out<=1;
   6962: out<=1;
   6963: out<=1;
   6964: out<=0;
   6965: out<=1;
   6966: out<=1;
   6967: out<=0;
   6968: out<=0;
   6969: out<=1;
   6970: out<=0;
   6971: out<=1;
   6972: out<=1;
   6973: out<=1;
   6974: out<=0;
   6975: out<=0;
   6976: out<=1;
   6977: out<=1;
   6978: out<=1;
   6979: out<=1;
   6980: out<=0;
   6981: out<=1;
   6982: out<=1;
   6983: out<=0;
   6984: out<=0;
   6985: out<=1;
   6986: out<=0;
   6987: out<=1;
   6988: out<=1;
   6989: out<=1;
   6990: out<=0;
   6991: out<=0;
   6992: out<=0;
   6993: out<=0;
   6994: out<=0;
   6995: out<=0;
   6996: out<=1;
   6997: out<=0;
   6998: out<=0;
   6999: out<=1;
   7000: out<=1;
   7001: out<=0;
   7002: out<=1;
   7003: out<=0;
   7004: out<=0;
   7005: out<=0;
   7006: out<=1;
   7007: out<=1;
   7008: out<=0;
   7009: out<=0;
   7010: out<=0;
   7011: out<=0;
   7012: out<=1;
   7013: out<=0;
   7014: out<=0;
   7015: out<=1;
   7016: out<=1;
   7017: out<=0;
   7018: out<=1;
   7019: out<=0;
   7020: out<=0;
   7021: out<=0;
   7022: out<=1;
   7023: out<=1;
   7024: out<=1;
   7025: out<=1;
   7026: out<=1;
   7027: out<=1;
   7028: out<=0;
   7029: out<=1;
   7030: out<=1;
   7031: out<=0;
   7032: out<=0;
   7033: out<=1;
   7034: out<=0;
   7035: out<=1;
   7036: out<=1;
   7037: out<=1;
   7038: out<=0;
   7039: out<=0;
   7040: out<=0;
   7041: out<=0;
   7042: out<=0;
   7043: out<=0;
   7044: out<=1;
   7045: out<=0;
   7046: out<=0;
   7047: out<=1;
   7048: out<=1;
   7049: out<=0;
   7050: out<=1;
   7051: out<=0;
   7052: out<=0;
   7053: out<=0;
   7054: out<=1;
   7055: out<=1;
   7056: out<=1;
   7057: out<=1;
   7058: out<=1;
   7059: out<=1;
   7060: out<=0;
   7061: out<=1;
   7062: out<=1;
   7063: out<=0;
   7064: out<=0;
   7065: out<=1;
   7066: out<=0;
   7067: out<=1;
   7068: out<=1;
   7069: out<=1;
   7070: out<=0;
   7071: out<=0;
   7072: out<=0;
   7073: out<=0;
   7074: out<=0;
   7075: out<=0;
   7076: out<=1;
   7077: out<=0;
   7078: out<=0;
   7079: out<=1;
   7080: out<=1;
   7081: out<=0;
   7082: out<=1;
   7083: out<=0;
   7084: out<=0;
   7085: out<=0;
   7086: out<=1;
   7087: out<=1;
   7088: out<=1;
   7089: out<=1;
   7090: out<=1;
   7091: out<=1;
   7092: out<=0;
   7093: out<=1;
   7094: out<=1;
   7095: out<=0;
   7096: out<=0;
   7097: out<=1;
   7098: out<=0;
   7099: out<=1;
   7100: out<=1;
   7101: out<=1;
   7102: out<=0;
   7103: out<=0;
   7104: out<=0;
   7105: out<=0;
   7106: out<=0;
   7107: out<=0;
   7108: out<=1;
   7109: out<=0;
   7110: out<=0;
   7111: out<=1;
   7112: out<=1;
   7113: out<=0;
   7114: out<=1;
   7115: out<=0;
   7116: out<=0;
   7117: out<=0;
   7118: out<=1;
   7119: out<=1;
   7120: out<=0;
   7121: out<=0;
   7122: out<=0;
   7123: out<=0;
   7124: out<=1;
   7125: out<=0;
   7126: out<=0;
   7127: out<=1;
   7128: out<=1;
   7129: out<=0;
   7130: out<=1;
   7131: out<=0;
   7132: out<=0;
   7133: out<=0;
   7134: out<=1;
   7135: out<=1;
   7136: out<=1;
   7137: out<=1;
   7138: out<=1;
   7139: out<=1;
   7140: out<=0;
   7141: out<=1;
   7142: out<=1;
   7143: out<=0;
   7144: out<=0;
   7145: out<=1;
   7146: out<=0;
   7147: out<=1;
   7148: out<=1;
   7149: out<=1;
   7150: out<=0;
   7151: out<=0;
   7152: out<=1;
   7153: out<=1;
   7154: out<=1;
   7155: out<=1;
   7156: out<=0;
   7157: out<=1;
   7158: out<=1;
   7159: out<=0;
   7160: out<=0;
   7161: out<=1;
   7162: out<=0;
   7163: out<=1;
   7164: out<=1;
   7165: out<=1;
   7166: out<=0;
   7167: out<=0;
   7168: out<=0;
   7169: out<=1;
   7170: out<=0;
   7171: out<=1;
   7172: out<=1;
   7173: out<=1;
   7174: out<=0;
   7175: out<=0;
   7176: out<=0;
   7177: out<=0;
   7178: out<=0;
   7179: out<=0;
   7180: out<=1;
   7181: out<=0;
   7182: out<=0;
   7183: out<=1;
   7184: out<=0;
   7185: out<=1;
   7186: out<=0;
   7187: out<=1;
   7188: out<=1;
   7189: out<=1;
   7190: out<=0;
   7191: out<=0;
   7192: out<=0;
   7193: out<=0;
   7194: out<=0;
   7195: out<=0;
   7196: out<=1;
   7197: out<=0;
   7198: out<=0;
   7199: out<=1;
   7200: out<=1;
   7201: out<=0;
   7202: out<=1;
   7203: out<=0;
   7204: out<=0;
   7205: out<=0;
   7206: out<=1;
   7207: out<=1;
   7208: out<=1;
   7209: out<=1;
   7210: out<=1;
   7211: out<=1;
   7212: out<=0;
   7213: out<=1;
   7214: out<=1;
   7215: out<=0;
   7216: out<=1;
   7217: out<=0;
   7218: out<=1;
   7219: out<=0;
   7220: out<=0;
   7221: out<=0;
   7222: out<=1;
   7223: out<=1;
   7224: out<=1;
   7225: out<=1;
   7226: out<=1;
   7227: out<=1;
   7228: out<=0;
   7229: out<=1;
   7230: out<=1;
   7231: out<=0;
   7232: out<=0;
   7233: out<=1;
   7234: out<=0;
   7235: out<=1;
   7236: out<=1;
   7237: out<=1;
   7238: out<=0;
   7239: out<=0;
   7240: out<=0;
   7241: out<=0;
   7242: out<=0;
   7243: out<=0;
   7244: out<=1;
   7245: out<=0;
   7246: out<=0;
   7247: out<=1;
   7248: out<=1;
   7249: out<=0;
   7250: out<=1;
   7251: out<=0;
   7252: out<=0;
   7253: out<=0;
   7254: out<=1;
   7255: out<=1;
   7256: out<=1;
   7257: out<=1;
   7258: out<=1;
   7259: out<=1;
   7260: out<=0;
   7261: out<=1;
   7262: out<=1;
   7263: out<=0;
   7264: out<=0;
   7265: out<=1;
   7266: out<=0;
   7267: out<=1;
   7268: out<=1;
   7269: out<=1;
   7270: out<=0;
   7271: out<=0;
   7272: out<=0;
   7273: out<=0;
   7274: out<=0;
   7275: out<=0;
   7276: out<=1;
   7277: out<=0;
   7278: out<=0;
   7279: out<=1;
   7280: out<=1;
   7281: out<=0;
   7282: out<=1;
   7283: out<=0;
   7284: out<=0;
   7285: out<=0;
   7286: out<=1;
   7287: out<=1;
   7288: out<=1;
   7289: out<=1;
   7290: out<=1;
   7291: out<=1;
   7292: out<=0;
   7293: out<=1;
   7294: out<=1;
   7295: out<=0;
   7296: out<=1;
   7297: out<=0;
   7298: out<=1;
   7299: out<=0;
   7300: out<=0;
   7301: out<=0;
   7302: out<=1;
   7303: out<=1;
   7304: out<=1;
   7305: out<=1;
   7306: out<=1;
   7307: out<=1;
   7308: out<=0;
   7309: out<=1;
   7310: out<=1;
   7311: out<=0;
   7312: out<=0;
   7313: out<=1;
   7314: out<=0;
   7315: out<=1;
   7316: out<=1;
   7317: out<=1;
   7318: out<=0;
   7319: out<=0;
   7320: out<=0;
   7321: out<=0;
   7322: out<=0;
   7323: out<=0;
   7324: out<=1;
   7325: out<=0;
   7326: out<=0;
   7327: out<=1;
   7328: out<=0;
   7329: out<=1;
   7330: out<=0;
   7331: out<=1;
   7332: out<=1;
   7333: out<=1;
   7334: out<=0;
   7335: out<=0;
   7336: out<=0;
   7337: out<=0;
   7338: out<=0;
   7339: out<=0;
   7340: out<=1;
   7341: out<=0;
   7342: out<=0;
   7343: out<=1;
   7344: out<=1;
   7345: out<=0;
   7346: out<=1;
   7347: out<=0;
   7348: out<=0;
   7349: out<=0;
   7350: out<=1;
   7351: out<=1;
   7352: out<=1;
   7353: out<=1;
   7354: out<=1;
   7355: out<=1;
   7356: out<=0;
   7357: out<=1;
   7358: out<=1;
   7359: out<=0;
   7360: out<=1;
   7361: out<=0;
   7362: out<=1;
   7363: out<=0;
   7364: out<=0;
   7365: out<=0;
   7366: out<=1;
   7367: out<=1;
   7368: out<=1;
   7369: out<=1;
   7370: out<=1;
   7371: out<=1;
   7372: out<=0;
   7373: out<=1;
   7374: out<=1;
   7375: out<=0;
   7376: out<=1;
   7377: out<=0;
   7378: out<=1;
   7379: out<=0;
   7380: out<=0;
   7381: out<=0;
   7382: out<=1;
   7383: out<=1;
   7384: out<=1;
   7385: out<=1;
   7386: out<=1;
   7387: out<=1;
   7388: out<=0;
   7389: out<=1;
   7390: out<=1;
   7391: out<=0;
   7392: out<=1;
   7393: out<=0;
   7394: out<=1;
   7395: out<=0;
   7396: out<=0;
   7397: out<=0;
   7398: out<=1;
   7399: out<=1;
   7400: out<=1;
   7401: out<=1;
   7402: out<=1;
   7403: out<=1;
   7404: out<=0;
   7405: out<=1;
   7406: out<=1;
   7407: out<=0;
   7408: out<=1;
   7409: out<=0;
   7410: out<=1;
   7411: out<=0;
   7412: out<=0;
   7413: out<=0;
   7414: out<=1;
   7415: out<=1;
   7416: out<=1;
   7417: out<=1;
   7418: out<=1;
   7419: out<=1;
   7420: out<=0;
   7421: out<=1;
   7422: out<=1;
   7423: out<=0;
   7424: out<=0;
   7425: out<=0;
   7426: out<=1;
   7427: out<=1;
   7428: out<=0;
   7429: out<=1;
   7430: out<=0;
   7431: out<=1;
   7432: out<=1;
   7433: out<=0;
   7434: out<=0;
   7435: out<=1;
   7436: out<=1;
   7437: out<=1;
   7438: out<=1;
   7439: out<=1;
   7440: out<=1;
   7441: out<=1;
   7442: out<=0;
   7443: out<=0;
   7444: out<=1;
   7445: out<=0;
   7446: out<=1;
   7447: out<=0;
   7448: out<=0;
   7449: out<=1;
   7450: out<=1;
   7451: out<=0;
   7452: out<=0;
   7453: out<=0;
   7454: out<=0;
   7455: out<=0;
   7456: out<=0;
   7457: out<=0;
   7458: out<=1;
   7459: out<=1;
   7460: out<=0;
   7461: out<=1;
   7462: out<=0;
   7463: out<=1;
   7464: out<=1;
   7465: out<=0;
   7466: out<=0;
   7467: out<=1;
   7468: out<=1;
   7469: out<=1;
   7470: out<=1;
   7471: out<=1;
   7472: out<=1;
   7473: out<=1;
   7474: out<=0;
   7475: out<=0;
   7476: out<=1;
   7477: out<=0;
   7478: out<=1;
   7479: out<=0;
   7480: out<=0;
   7481: out<=1;
   7482: out<=1;
   7483: out<=0;
   7484: out<=0;
   7485: out<=0;
   7486: out<=0;
   7487: out<=0;
   7488: out<=0;
   7489: out<=0;
   7490: out<=1;
   7491: out<=1;
   7492: out<=0;
   7493: out<=1;
   7494: out<=0;
   7495: out<=1;
   7496: out<=1;
   7497: out<=0;
   7498: out<=0;
   7499: out<=1;
   7500: out<=1;
   7501: out<=1;
   7502: out<=1;
   7503: out<=1;
   7504: out<=0;
   7505: out<=0;
   7506: out<=1;
   7507: out<=1;
   7508: out<=0;
   7509: out<=1;
   7510: out<=0;
   7511: out<=1;
   7512: out<=1;
   7513: out<=0;
   7514: out<=0;
   7515: out<=1;
   7516: out<=1;
   7517: out<=1;
   7518: out<=1;
   7519: out<=1;
   7520: out<=1;
   7521: out<=1;
   7522: out<=0;
   7523: out<=0;
   7524: out<=1;
   7525: out<=0;
   7526: out<=1;
   7527: out<=0;
   7528: out<=0;
   7529: out<=1;
   7530: out<=1;
   7531: out<=0;
   7532: out<=0;
   7533: out<=0;
   7534: out<=0;
   7535: out<=0;
   7536: out<=1;
   7537: out<=1;
   7538: out<=0;
   7539: out<=0;
   7540: out<=1;
   7541: out<=0;
   7542: out<=1;
   7543: out<=0;
   7544: out<=0;
   7545: out<=1;
   7546: out<=1;
   7547: out<=0;
   7548: out<=0;
   7549: out<=0;
   7550: out<=0;
   7551: out<=0;
   7552: out<=1;
   7553: out<=1;
   7554: out<=0;
   7555: out<=0;
   7556: out<=1;
   7557: out<=0;
   7558: out<=1;
   7559: out<=0;
   7560: out<=0;
   7561: out<=1;
   7562: out<=1;
   7563: out<=0;
   7564: out<=0;
   7565: out<=0;
   7566: out<=0;
   7567: out<=0;
   7568: out<=1;
   7569: out<=1;
   7570: out<=0;
   7571: out<=0;
   7572: out<=1;
   7573: out<=0;
   7574: out<=1;
   7575: out<=0;
   7576: out<=0;
   7577: out<=1;
   7578: out<=1;
   7579: out<=0;
   7580: out<=0;
   7581: out<=0;
   7582: out<=0;
   7583: out<=0;
   7584: out<=1;
   7585: out<=1;
   7586: out<=0;
   7587: out<=0;
   7588: out<=1;
   7589: out<=0;
   7590: out<=1;
   7591: out<=0;
   7592: out<=0;
   7593: out<=1;
   7594: out<=1;
   7595: out<=0;
   7596: out<=0;
   7597: out<=0;
   7598: out<=0;
   7599: out<=0;
   7600: out<=1;
   7601: out<=1;
   7602: out<=0;
   7603: out<=0;
   7604: out<=1;
   7605: out<=0;
   7606: out<=1;
   7607: out<=0;
   7608: out<=0;
   7609: out<=1;
   7610: out<=1;
   7611: out<=0;
   7612: out<=0;
   7613: out<=0;
   7614: out<=0;
   7615: out<=0;
   7616: out<=1;
   7617: out<=1;
   7618: out<=0;
   7619: out<=0;
   7620: out<=1;
   7621: out<=0;
   7622: out<=1;
   7623: out<=0;
   7624: out<=0;
   7625: out<=1;
   7626: out<=1;
   7627: out<=0;
   7628: out<=0;
   7629: out<=0;
   7630: out<=0;
   7631: out<=0;
   7632: out<=0;
   7633: out<=0;
   7634: out<=1;
   7635: out<=1;
   7636: out<=0;
   7637: out<=1;
   7638: out<=0;
   7639: out<=1;
   7640: out<=1;
   7641: out<=0;
   7642: out<=0;
   7643: out<=1;
   7644: out<=1;
   7645: out<=1;
   7646: out<=1;
   7647: out<=1;
   7648: out<=0;
   7649: out<=0;
   7650: out<=1;
   7651: out<=1;
   7652: out<=0;
   7653: out<=1;
   7654: out<=0;
   7655: out<=1;
   7656: out<=1;
   7657: out<=0;
   7658: out<=0;
   7659: out<=1;
   7660: out<=1;
   7661: out<=1;
   7662: out<=1;
   7663: out<=1;
   7664: out<=1;
   7665: out<=1;
   7666: out<=0;
   7667: out<=0;
   7668: out<=1;
   7669: out<=0;
   7670: out<=1;
   7671: out<=0;
   7672: out<=0;
   7673: out<=1;
   7674: out<=1;
   7675: out<=0;
   7676: out<=0;
   7677: out<=0;
   7678: out<=0;
   7679: out<=0;
   7680: out<=1;
   7681: out<=1;
   7682: out<=1;
   7683: out<=1;
   7684: out<=1;
   7685: out<=0;
   7686: out<=0;
   7687: out<=1;
   7688: out<=1;
   7689: out<=0;
   7690: out<=1;
   7691: out<=0;
   7692: out<=1;
   7693: out<=1;
   7694: out<=0;
   7695: out<=0;
   7696: out<=0;
   7697: out<=0;
   7698: out<=0;
   7699: out<=0;
   7700: out<=0;
   7701: out<=1;
   7702: out<=1;
   7703: out<=0;
   7704: out<=0;
   7705: out<=1;
   7706: out<=0;
   7707: out<=1;
   7708: out<=0;
   7709: out<=0;
   7710: out<=1;
   7711: out<=1;
   7712: out<=0;
   7713: out<=0;
   7714: out<=0;
   7715: out<=0;
   7716: out<=0;
   7717: out<=1;
   7718: out<=1;
   7719: out<=0;
   7720: out<=0;
   7721: out<=1;
   7722: out<=0;
   7723: out<=1;
   7724: out<=0;
   7725: out<=0;
   7726: out<=1;
   7727: out<=1;
   7728: out<=1;
   7729: out<=1;
   7730: out<=1;
   7731: out<=1;
   7732: out<=1;
   7733: out<=0;
   7734: out<=0;
   7735: out<=1;
   7736: out<=1;
   7737: out<=0;
   7738: out<=1;
   7739: out<=0;
   7740: out<=1;
   7741: out<=1;
   7742: out<=0;
   7743: out<=0;
   7744: out<=1;
   7745: out<=1;
   7746: out<=1;
   7747: out<=1;
   7748: out<=1;
   7749: out<=0;
   7750: out<=0;
   7751: out<=1;
   7752: out<=1;
   7753: out<=0;
   7754: out<=1;
   7755: out<=0;
   7756: out<=1;
   7757: out<=1;
   7758: out<=0;
   7759: out<=0;
   7760: out<=1;
   7761: out<=1;
   7762: out<=1;
   7763: out<=1;
   7764: out<=1;
   7765: out<=0;
   7766: out<=0;
   7767: out<=1;
   7768: out<=1;
   7769: out<=0;
   7770: out<=1;
   7771: out<=0;
   7772: out<=1;
   7773: out<=1;
   7774: out<=0;
   7775: out<=0;
   7776: out<=1;
   7777: out<=1;
   7778: out<=1;
   7779: out<=1;
   7780: out<=1;
   7781: out<=0;
   7782: out<=0;
   7783: out<=1;
   7784: out<=1;
   7785: out<=0;
   7786: out<=1;
   7787: out<=0;
   7788: out<=1;
   7789: out<=1;
   7790: out<=0;
   7791: out<=0;
   7792: out<=1;
   7793: out<=1;
   7794: out<=1;
   7795: out<=1;
   7796: out<=1;
   7797: out<=0;
   7798: out<=0;
   7799: out<=1;
   7800: out<=1;
   7801: out<=0;
   7802: out<=1;
   7803: out<=0;
   7804: out<=1;
   7805: out<=1;
   7806: out<=0;
   7807: out<=0;
   7808: out<=0;
   7809: out<=0;
   7810: out<=0;
   7811: out<=0;
   7812: out<=0;
   7813: out<=1;
   7814: out<=1;
   7815: out<=0;
   7816: out<=0;
   7817: out<=1;
   7818: out<=0;
   7819: out<=1;
   7820: out<=0;
   7821: out<=0;
   7822: out<=1;
   7823: out<=1;
   7824: out<=0;
   7825: out<=0;
   7826: out<=0;
   7827: out<=0;
   7828: out<=0;
   7829: out<=1;
   7830: out<=1;
   7831: out<=0;
   7832: out<=0;
   7833: out<=1;
   7834: out<=0;
   7835: out<=1;
   7836: out<=0;
   7837: out<=0;
   7838: out<=1;
   7839: out<=1;
   7840: out<=1;
   7841: out<=1;
   7842: out<=1;
   7843: out<=1;
   7844: out<=1;
   7845: out<=0;
   7846: out<=0;
   7847: out<=1;
   7848: out<=1;
   7849: out<=0;
   7850: out<=1;
   7851: out<=0;
   7852: out<=1;
   7853: out<=1;
   7854: out<=0;
   7855: out<=0;
   7856: out<=1;
   7857: out<=1;
   7858: out<=1;
   7859: out<=1;
   7860: out<=1;
   7861: out<=0;
   7862: out<=0;
   7863: out<=1;
   7864: out<=1;
   7865: out<=0;
   7866: out<=1;
   7867: out<=0;
   7868: out<=1;
   7869: out<=1;
   7870: out<=0;
   7871: out<=0;
   7872: out<=0;
   7873: out<=0;
   7874: out<=0;
   7875: out<=0;
   7876: out<=0;
   7877: out<=1;
   7878: out<=1;
   7879: out<=0;
   7880: out<=0;
   7881: out<=1;
   7882: out<=0;
   7883: out<=1;
   7884: out<=0;
   7885: out<=0;
   7886: out<=1;
   7887: out<=1;
   7888: out<=1;
   7889: out<=1;
   7890: out<=1;
   7891: out<=1;
   7892: out<=1;
   7893: out<=0;
   7894: out<=0;
   7895: out<=1;
   7896: out<=1;
   7897: out<=0;
   7898: out<=1;
   7899: out<=0;
   7900: out<=1;
   7901: out<=1;
   7902: out<=0;
   7903: out<=0;
   7904: out<=0;
   7905: out<=0;
   7906: out<=0;
   7907: out<=0;
   7908: out<=0;
   7909: out<=1;
   7910: out<=1;
   7911: out<=0;
   7912: out<=0;
   7913: out<=1;
   7914: out<=0;
   7915: out<=1;
   7916: out<=0;
   7917: out<=0;
   7918: out<=1;
   7919: out<=1;
   7920: out<=1;
   7921: out<=1;
   7922: out<=1;
   7923: out<=1;
   7924: out<=1;
   7925: out<=0;
   7926: out<=0;
   7927: out<=1;
   7928: out<=1;
   7929: out<=0;
   7930: out<=1;
   7931: out<=0;
   7932: out<=1;
   7933: out<=1;
   7934: out<=0;
   7935: out<=0;
   7936: out<=1;
   7937: out<=0;
   7938: out<=0;
   7939: out<=1;
   7940: out<=0;
   7941: out<=0;
   7942: out<=0;
   7943: out<=0;
   7944: out<=0;
   7945: out<=0;
   7946: out<=1;
   7947: out<=1;
   7948: out<=1;
   7949: out<=0;
   7950: out<=1;
   7951: out<=0;
   7952: out<=1;
   7953: out<=0;
   7954: out<=0;
   7955: out<=1;
   7956: out<=0;
   7957: out<=0;
   7958: out<=0;
   7959: out<=0;
   7960: out<=0;
   7961: out<=0;
   7962: out<=1;
   7963: out<=1;
   7964: out<=1;
   7965: out<=0;
   7966: out<=1;
   7967: out<=0;
   7968: out<=1;
   7969: out<=0;
   7970: out<=0;
   7971: out<=1;
   7972: out<=0;
   7973: out<=0;
   7974: out<=0;
   7975: out<=0;
   7976: out<=0;
   7977: out<=0;
   7978: out<=1;
   7979: out<=1;
   7980: out<=1;
   7981: out<=0;
   7982: out<=1;
   7983: out<=0;
   7984: out<=1;
   7985: out<=0;
   7986: out<=0;
   7987: out<=1;
   7988: out<=0;
   7989: out<=0;
   7990: out<=0;
   7991: out<=0;
   7992: out<=0;
   7993: out<=0;
   7994: out<=1;
   7995: out<=1;
   7996: out<=1;
   7997: out<=0;
   7998: out<=1;
   7999: out<=0;
   8000: out<=1;
   8001: out<=0;
   8002: out<=0;
   8003: out<=1;
   8004: out<=0;
   8005: out<=0;
   8006: out<=0;
   8007: out<=0;
   8008: out<=0;
   8009: out<=0;
   8010: out<=1;
   8011: out<=1;
   8012: out<=1;
   8013: out<=0;
   8014: out<=1;
   8015: out<=0;
   8016: out<=0;
   8017: out<=1;
   8018: out<=1;
   8019: out<=0;
   8020: out<=1;
   8021: out<=1;
   8022: out<=1;
   8023: out<=1;
   8024: out<=1;
   8025: out<=1;
   8026: out<=0;
   8027: out<=0;
   8028: out<=0;
   8029: out<=1;
   8030: out<=0;
   8031: out<=1;
   8032: out<=0;
   8033: out<=1;
   8034: out<=1;
   8035: out<=0;
   8036: out<=1;
   8037: out<=1;
   8038: out<=1;
   8039: out<=1;
   8040: out<=1;
   8041: out<=1;
   8042: out<=0;
   8043: out<=0;
   8044: out<=0;
   8045: out<=1;
   8046: out<=0;
   8047: out<=1;
   8048: out<=1;
   8049: out<=0;
   8050: out<=0;
   8051: out<=1;
   8052: out<=0;
   8053: out<=0;
   8054: out<=0;
   8055: out<=0;
   8056: out<=0;
   8057: out<=0;
   8058: out<=1;
   8059: out<=1;
   8060: out<=1;
   8061: out<=0;
   8062: out<=1;
   8063: out<=0;
   8064: out<=0;
   8065: out<=1;
   8066: out<=1;
   8067: out<=0;
   8068: out<=1;
   8069: out<=1;
   8070: out<=1;
   8071: out<=1;
   8072: out<=1;
   8073: out<=1;
   8074: out<=0;
   8075: out<=0;
   8076: out<=0;
   8077: out<=1;
   8078: out<=0;
   8079: out<=1;
   8080: out<=1;
   8081: out<=0;
   8082: out<=0;
   8083: out<=1;
   8084: out<=0;
   8085: out<=0;
   8086: out<=0;
   8087: out<=0;
   8088: out<=0;
   8089: out<=0;
   8090: out<=1;
   8091: out<=1;
   8092: out<=1;
   8093: out<=0;
   8094: out<=1;
   8095: out<=0;
   8096: out<=0;
   8097: out<=1;
   8098: out<=1;
   8099: out<=0;
   8100: out<=1;
   8101: out<=1;
   8102: out<=1;
   8103: out<=1;
   8104: out<=1;
   8105: out<=1;
   8106: out<=0;
   8107: out<=0;
   8108: out<=0;
   8109: out<=1;
   8110: out<=0;
   8111: out<=1;
   8112: out<=1;
   8113: out<=0;
   8114: out<=0;
   8115: out<=1;
   8116: out<=0;
   8117: out<=0;
   8118: out<=0;
   8119: out<=0;
   8120: out<=0;
   8121: out<=0;
   8122: out<=1;
   8123: out<=1;
   8124: out<=1;
   8125: out<=0;
   8126: out<=1;
   8127: out<=0;
   8128: out<=0;
   8129: out<=1;
   8130: out<=1;
   8131: out<=0;
   8132: out<=1;
   8133: out<=1;
   8134: out<=1;
   8135: out<=1;
   8136: out<=1;
   8137: out<=1;
   8138: out<=0;
   8139: out<=0;
   8140: out<=0;
   8141: out<=1;
   8142: out<=0;
   8143: out<=1;
   8144: out<=0;
   8145: out<=1;
   8146: out<=1;
   8147: out<=0;
   8148: out<=1;
   8149: out<=1;
   8150: out<=1;
   8151: out<=1;
   8152: out<=1;
   8153: out<=1;
   8154: out<=0;
   8155: out<=0;
   8156: out<=0;
   8157: out<=1;
   8158: out<=0;
   8159: out<=1;
   8160: out<=1;
   8161: out<=0;
   8162: out<=0;
   8163: out<=1;
   8164: out<=0;
   8165: out<=0;
   8166: out<=0;
   8167: out<=0;
   8168: out<=0;
   8169: out<=0;
   8170: out<=1;
   8171: out<=1;
   8172: out<=1;
   8173: out<=0;
   8174: out<=1;
   8175: out<=0;
   8176: out<=1;
   8177: out<=0;
   8178: out<=0;
   8179: out<=1;
   8180: out<=0;
   8181: out<=0;
   8182: out<=0;
   8183: out<=0;
   8184: out<=0;
   8185: out<=0;
   8186: out<=1;
   8187: out<=1;
   8188: out<=1;
   8189: out<=0;
   8190: out<=1;
   8191: out<=0;
   8192: out<=0;
   8193: out<=1;
   8194: out<=0;
   8195: out<=1;
   8196: out<=1;
   8197: out<=1;
   8198: out<=0;
   8199: out<=0;
   8200: out<=0;
   8201: out<=0;
   8202: out<=0;
   8203: out<=0;
   8204: out<=1;
   8205: out<=0;
   8206: out<=0;
   8207: out<=1;
   8208: out<=0;
   8209: out<=1;
   8210: out<=0;
   8211: out<=1;
   8212: out<=1;
   8213: out<=1;
   8214: out<=0;
   8215: out<=0;
   8216: out<=0;
   8217: out<=0;
   8218: out<=0;
   8219: out<=0;
   8220: out<=1;
   8221: out<=0;
   8222: out<=0;
   8223: out<=1;
   8224: out<=0;
   8225: out<=1;
   8226: out<=0;
   8227: out<=1;
   8228: out<=1;
   8229: out<=1;
   8230: out<=0;
   8231: out<=0;
   8232: out<=0;
   8233: out<=0;
   8234: out<=0;
   8235: out<=0;
   8236: out<=1;
   8237: out<=0;
   8238: out<=0;
   8239: out<=1;
   8240: out<=0;
   8241: out<=1;
   8242: out<=0;
   8243: out<=1;
   8244: out<=1;
   8245: out<=1;
   8246: out<=0;
   8247: out<=0;
   8248: out<=0;
   8249: out<=0;
   8250: out<=0;
   8251: out<=0;
   8252: out<=1;
   8253: out<=0;
   8254: out<=0;
   8255: out<=1;
   8256: out<=0;
   8257: out<=1;
   8258: out<=0;
   8259: out<=1;
   8260: out<=1;
   8261: out<=1;
   8262: out<=0;
   8263: out<=0;
   8264: out<=0;
   8265: out<=0;
   8266: out<=0;
   8267: out<=0;
   8268: out<=1;
   8269: out<=0;
   8270: out<=0;
   8271: out<=1;
   8272: out<=1;
   8273: out<=0;
   8274: out<=1;
   8275: out<=0;
   8276: out<=0;
   8277: out<=0;
   8278: out<=1;
   8279: out<=1;
   8280: out<=1;
   8281: out<=1;
   8282: out<=1;
   8283: out<=1;
   8284: out<=0;
   8285: out<=1;
   8286: out<=1;
   8287: out<=0;
   8288: out<=1;
   8289: out<=0;
   8290: out<=1;
   8291: out<=0;
   8292: out<=0;
   8293: out<=0;
   8294: out<=1;
   8295: out<=1;
   8296: out<=1;
   8297: out<=1;
   8298: out<=1;
   8299: out<=1;
   8300: out<=0;
   8301: out<=1;
   8302: out<=1;
   8303: out<=0;
   8304: out<=0;
   8305: out<=1;
   8306: out<=0;
   8307: out<=1;
   8308: out<=1;
   8309: out<=1;
   8310: out<=0;
   8311: out<=0;
   8312: out<=0;
   8313: out<=0;
   8314: out<=0;
   8315: out<=0;
   8316: out<=1;
   8317: out<=0;
   8318: out<=0;
   8319: out<=1;
   8320: out<=0;
   8321: out<=1;
   8322: out<=0;
   8323: out<=1;
   8324: out<=1;
   8325: out<=1;
   8326: out<=0;
   8327: out<=0;
   8328: out<=0;
   8329: out<=0;
   8330: out<=0;
   8331: out<=0;
   8332: out<=1;
   8333: out<=0;
   8334: out<=0;
   8335: out<=1;
   8336: out<=1;
   8337: out<=0;
   8338: out<=1;
   8339: out<=0;
   8340: out<=0;
   8341: out<=0;
   8342: out<=1;
   8343: out<=1;
   8344: out<=1;
   8345: out<=1;
   8346: out<=1;
   8347: out<=1;
   8348: out<=0;
   8349: out<=1;
   8350: out<=1;
   8351: out<=0;
   8352: out<=0;
   8353: out<=1;
   8354: out<=0;
   8355: out<=1;
   8356: out<=1;
   8357: out<=1;
   8358: out<=0;
   8359: out<=0;
   8360: out<=0;
   8361: out<=0;
   8362: out<=0;
   8363: out<=0;
   8364: out<=1;
   8365: out<=0;
   8366: out<=0;
   8367: out<=1;
   8368: out<=1;
   8369: out<=0;
   8370: out<=1;
   8371: out<=0;
   8372: out<=0;
   8373: out<=0;
   8374: out<=1;
   8375: out<=1;
   8376: out<=1;
   8377: out<=1;
   8378: out<=1;
   8379: out<=1;
   8380: out<=0;
   8381: out<=1;
   8382: out<=1;
   8383: out<=0;
   8384: out<=0;
   8385: out<=1;
   8386: out<=0;
   8387: out<=1;
   8388: out<=1;
   8389: out<=1;
   8390: out<=0;
   8391: out<=0;
   8392: out<=0;
   8393: out<=0;
   8394: out<=0;
   8395: out<=0;
   8396: out<=1;
   8397: out<=0;
   8398: out<=0;
   8399: out<=1;
   8400: out<=0;
   8401: out<=1;
   8402: out<=0;
   8403: out<=1;
   8404: out<=1;
   8405: out<=1;
   8406: out<=0;
   8407: out<=0;
   8408: out<=0;
   8409: out<=0;
   8410: out<=0;
   8411: out<=0;
   8412: out<=1;
   8413: out<=0;
   8414: out<=0;
   8415: out<=1;
   8416: out<=1;
   8417: out<=0;
   8418: out<=1;
   8419: out<=0;
   8420: out<=0;
   8421: out<=0;
   8422: out<=1;
   8423: out<=1;
   8424: out<=1;
   8425: out<=1;
   8426: out<=1;
   8427: out<=1;
   8428: out<=0;
   8429: out<=1;
   8430: out<=1;
   8431: out<=0;
   8432: out<=1;
   8433: out<=0;
   8434: out<=1;
   8435: out<=0;
   8436: out<=0;
   8437: out<=0;
   8438: out<=1;
   8439: out<=1;
   8440: out<=1;
   8441: out<=1;
   8442: out<=1;
   8443: out<=1;
   8444: out<=0;
   8445: out<=1;
   8446: out<=1;
   8447: out<=0;
   8448: out<=0;
   8449: out<=0;
   8450: out<=1;
   8451: out<=1;
   8452: out<=0;
   8453: out<=1;
   8454: out<=0;
   8455: out<=1;
   8456: out<=1;
   8457: out<=0;
   8458: out<=0;
   8459: out<=1;
   8460: out<=1;
   8461: out<=1;
   8462: out<=1;
   8463: out<=1;
   8464: out<=1;
   8465: out<=1;
   8466: out<=0;
   8467: out<=0;
   8468: out<=1;
   8469: out<=0;
   8470: out<=1;
   8471: out<=0;
   8472: out<=0;
   8473: out<=1;
   8474: out<=1;
   8475: out<=0;
   8476: out<=0;
   8477: out<=0;
   8478: out<=0;
   8479: out<=0;
   8480: out<=1;
   8481: out<=1;
   8482: out<=0;
   8483: out<=0;
   8484: out<=1;
   8485: out<=0;
   8486: out<=1;
   8487: out<=0;
   8488: out<=0;
   8489: out<=1;
   8490: out<=1;
   8491: out<=0;
   8492: out<=0;
   8493: out<=0;
   8494: out<=0;
   8495: out<=0;
   8496: out<=0;
   8497: out<=0;
   8498: out<=1;
   8499: out<=1;
   8500: out<=0;
   8501: out<=1;
   8502: out<=0;
   8503: out<=1;
   8504: out<=1;
   8505: out<=0;
   8506: out<=0;
   8507: out<=1;
   8508: out<=1;
   8509: out<=1;
   8510: out<=1;
   8511: out<=1;
   8512: out<=0;
   8513: out<=0;
   8514: out<=1;
   8515: out<=1;
   8516: out<=0;
   8517: out<=1;
   8518: out<=0;
   8519: out<=1;
   8520: out<=1;
   8521: out<=0;
   8522: out<=0;
   8523: out<=1;
   8524: out<=1;
   8525: out<=1;
   8526: out<=1;
   8527: out<=1;
   8528: out<=0;
   8529: out<=0;
   8530: out<=1;
   8531: out<=1;
   8532: out<=0;
   8533: out<=1;
   8534: out<=0;
   8535: out<=1;
   8536: out<=1;
   8537: out<=0;
   8538: out<=0;
   8539: out<=1;
   8540: out<=1;
   8541: out<=1;
   8542: out<=1;
   8543: out<=1;
   8544: out<=0;
   8545: out<=0;
   8546: out<=1;
   8547: out<=1;
   8548: out<=0;
   8549: out<=1;
   8550: out<=0;
   8551: out<=1;
   8552: out<=1;
   8553: out<=0;
   8554: out<=0;
   8555: out<=1;
   8556: out<=1;
   8557: out<=1;
   8558: out<=1;
   8559: out<=1;
   8560: out<=0;
   8561: out<=0;
   8562: out<=1;
   8563: out<=1;
   8564: out<=0;
   8565: out<=1;
   8566: out<=0;
   8567: out<=1;
   8568: out<=1;
   8569: out<=0;
   8570: out<=0;
   8571: out<=1;
   8572: out<=1;
   8573: out<=1;
   8574: out<=1;
   8575: out<=1;
   8576: out<=0;
   8577: out<=0;
   8578: out<=1;
   8579: out<=1;
   8580: out<=0;
   8581: out<=1;
   8582: out<=0;
   8583: out<=1;
   8584: out<=1;
   8585: out<=0;
   8586: out<=0;
   8587: out<=1;
   8588: out<=1;
   8589: out<=1;
   8590: out<=1;
   8591: out<=1;
   8592: out<=0;
   8593: out<=0;
   8594: out<=1;
   8595: out<=1;
   8596: out<=0;
   8597: out<=1;
   8598: out<=0;
   8599: out<=1;
   8600: out<=1;
   8601: out<=0;
   8602: out<=0;
   8603: out<=1;
   8604: out<=1;
   8605: out<=1;
   8606: out<=1;
   8607: out<=1;
   8608: out<=1;
   8609: out<=1;
   8610: out<=0;
   8611: out<=0;
   8612: out<=1;
   8613: out<=0;
   8614: out<=1;
   8615: out<=0;
   8616: out<=0;
   8617: out<=1;
   8618: out<=1;
   8619: out<=0;
   8620: out<=0;
   8621: out<=0;
   8622: out<=0;
   8623: out<=0;
   8624: out<=1;
   8625: out<=1;
   8626: out<=0;
   8627: out<=0;
   8628: out<=1;
   8629: out<=0;
   8630: out<=1;
   8631: out<=0;
   8632: out<=0;
   8633: out<=1;
   8634: out<=1;
   8635: out<=0;
   8636: out<=0;
   8637: out<=0;
   8638: out<=0;
   8639: out<=0;
   8640: out<=0;
   8641: out<=0;
   8642: out<=1;
   8643: out<=1;
   8644: out<=0;
   8645: out<=1;
   8646: out<=0;
   8647: out<=1;
   8648: out<=1;
   8649: out<=0;
   8650: out<=0;
   8651: out<=1;
   8652: out<=1;
   8653: out<=1;
   8654: out<=1;
   8655: out<=1;
   8656: out<=1;
   8657: out<=1;
   8658: out<=0;
   8659: out<=0;
   8660: out<=1;
   8661: out<=0;
   8662: out<=1;
   8663: out<=0;
   8664: out<=0;
   8665: out<=1;
   8666: out<=1;
   8667: out<=0;
   8668: out<=0;
   8669: out<=0;
   8670: out<=0;
   8671: out<=0;
   8672: out<=0;
   8673: out<=0;
   8674: out<=1;
   8675: out<=1;
   8676: out<=0;
   8677: out<=1;
   8678: out<=0;
   8679: out<=1;
   8680: out<=1;
   8681: out<=0;
   8682: out<=0;
   8683: out<=1;
   8684: out<=1;
   8685: out<=1;
   8686: out<=1;
   8687: out<=1;
   8688: out<=1;
   8689: out<=1;
   8690: out<=0;
   8691: out<=0;
   8692: out<=1;
   8693: out<=0;
   8694: out<=1;
   8695: out<=0;
   8696: out<=0;
   8697: out<=1;
   8698: out<=1;
   8699: out<=0;
   8700: out<=0;
   8701: out<=0;
   8702: out<=0;
   8703: out<=0;
   8704: out<=0;
   8705: out<=0;
   8706: out<=0;
   8707: out<=0;
   8708: out<=0;
   8709: out<=1;
   8710: out<=1;
   8711: out<=0;
   8712: out<=0;
   8713: out<=1;
   8714: out<=0;
   8715: out<=1;
   8716: out<=0;
   8717: out<=0;
   8718: out<=1;
   8719: out<=1;
   8720: out<=1;
   8721: out<=1;
   8722: out<=1;
   8723: out<=1;
   8724: out<=1;
   8725: out<=0;
   8726: out<=0;
   8727: out<=1;
   8728: out<=1;
   8729: out<=0;
   8730: out<=1;
   8731: out<=0;
   8732: out<=1;
   8733: out<=1;
   8734: out<=0;
   8735: out<=0;
   8736: out<=0;
   8737: out<=0;
   8738: out<=0;
   8739: out<=0;
   8740: out<=0;
   8741: out<=1;
   8742: out<=1;
   8743: out<=0;
   8744: out<=0;
   8745: out<=1;
   8746: out<=0;
   8747: out<=1;
   8748: out<=0;
   8749: out<=0;
   8750: out<=1;
   8751: out<=1;
   8752: out<=1;
   8753: out<=1;
   8754: out<=1;
   8755: out<=1;
   8756: out<=1;
   8757: out<=0;
   8758: out<=0;
   8759: out<=1;
   8760: out<=1;
   8761: out<=0;
   8762: out<=1;
   8763: out<=0;
   8764: out<=1;
   8765: out<=1;
   8766: out<=0;
   8767: out<=0;
   8768: out<=0;
   8769: out<=0;
   8770: out<=0;
   8771: out<=0;
   8772: out<=0;
   8773: out<=1;
   8774: out<=1;
   8775: out<=0;
   8776: out<=0;
   8777: out<=1;
   8778: out<=0;
   8779: out<=1;
   8780: out<=0;
   8781: out<=0;
   8782: out<=1;
   8783: out<=1;
   8784: out<=0;
   8785: out<=0;
   8786: out<=0;
   8787: out<=0;
   8788: out<=0;
   8789: out<=1;
   8790: out<=1;
   8791: out<=0;
   8792: out<=0;
   8793: out<=1;
   8794: out<=0;
   8795: out<=1;
   8796: out<=0;
   8797: out<=0;
   8798: out<=1;
   8799: out<=1;
   8800: out<=1;
   8801: out<=1;
   8802: out<=1;
   8803: out<=1;
   8804: out<=1;
   8805: out<=0;
   8806: out<=0;
   8807: out<=1;
   8808: out<=1;
   8809: out<=0;
   8810: out<=1;
   8811: out<=0;
   8812: out<=1;
   8813: out<=1;
   8814: out<=0;
   8815: out<=0;
   8816: out<=1;
   8817: out<=1;
   8818: out<=1;
   8819: out<=1;
   8820: out<=1;
   8821: out<=0;
   8822: out<=0;
   8823: out<=1;
   8824: out<=1;
   8825: out<=0;
   8826: out<=1;
   8827: out<=0;
   8828: out<=1;
   8829: out<=1;
   8830: out<=0;
   8831: out<=0;
   8832: out<=0;
   8833: out<=0;
   8834: out<=0;
   8835: out<=0;
   8836: out<=0;
   8837: out<=1;
   8838: out<=1;
   8839: out<=0;
   8840: out<=0;
   8841: out<=1;
   8842: out<=0;
   8843: out<=1;
   8844: out<=0;
   8845: out<=0;
   8846: out<=1;
   8847: out<=1;
   8848: out<=0;
   8849: out<=0;
   8850: out<=0;
   8851: out<=0;
   8852: out<=0;
   8853: out<=1;
   8854: out<=1;
   8855: out<=0;
   8856: out<=0;
   8857: out<=1;
   8858: out<=0;
   8859: out<=1;
   8860: out<=0;
   8861: out<=0;
   8862: out<=1;
   8863: out<=1;
   8864: out<=0;
   8865: out<=0;
   8866: out<=0;
   8867: out<=0;
   8868: out<=0;
   8869: out<=1;
   8870: out<=1;
   8871: out<=0;
   8872: out<=0;
   8873: out<=1;
   8874: out<=0;
   8875: out<=1;
   8876: out<=0;
   8877: out<=0;
   8878: out<=1;
   8879: out<=1;
   8880: out<=0;
   8881: out<=0;
   8882: out<=0;
   8883: out<=0;
   8884: out<=0;
   8885: out<=1;
   8886: out<=1;
   8887: out<=0;
   8888: out<=0;
   8889: out<=1;
   8890: out<=0;
   8891: out<=1;
   8892: out<=0;
   8893: out<=0;
   8894: out<=1;
   8895: out<=1;
   8896: out<=0;
   8897: out<=0;
   8898: out<=0;
   8899: out<=0;
   8900: out<=0;
   8901: out<=1;
   8902: out<=1;
   8903: out<=0;
   8904: out<=0;
   8905: out<=1;
   8906: out<=0;
   8907: out<=1;
   8908: out<=0;
   8909: out<=0;
   8910: out<=1;
   8911: out<=1;
   8912: out<=1;
   8913: out<=1;
   8914: out<=1;
   8915: out<=1;
   8916: out<=1;
   8917: out<=0;
   8918: out<=0;
   8919: out<=1;
   8920: out<=1;
   8921: out<=0;
   8922: out<=1;
   8923: out<=0;
   8924: out<=1;
   8925: out<=1;
   8926: out<=0;
   8927: out<=0;
   8928: out<=1;
   8929: out<=1;
   8930: out<=1;
   8931: out<=1;
   8932: out<=1;
   8933: out<=0;
   8934: out<=0;
   8935: out<=1;
   8936: out<=1;
   8937: out<=0;
   8938: out<=1;
   8939: out<=0;
   8940: out<=1;
   8941: out<=1;
   8942: out<=0;
   8943: out<=0;
   8944: out<=0;
   8945: out<=0;
   8946: out<=0;
   8947: out<=0;
   8948: out<=0;
   8949: out<=1;
   8950: out<=1;
   8951: out<=0;
   8952: out<=0;
   8953: out<=1;
   8954: out<=0;
   8955: out<=1;
   8956: out<=0;
   8957: out<=0;
   8958: out<=1;
   8959: out<=1;
   8960: out<=0;
   8961: out<=1;
   8962: out<=1;
   8963: out<=0;
   8964: out<=1;
   8965: out<=1;
   8966: out<=1;
   8967: out<=1;
   8968: out<=1;
   8969: out<=1;
   8970: out<=0;
   8971: out<=0;
   8972: out<=0;
   8973: out<=1;
   8974: out<=0;
   8975: out<=1;
   8976: out<=0;
   8977: out<=1;
   8978: out<=1;
   8979: out<=0;
   8980: out<=1;
   8981: out<=1;
   8982: out<=1;
   8983: out<=1;
   8984: out<=1;
   8985: out<=1;
   8986: out<=0;
   8987: out<=0;
   8988: out<=0;
   8989: out<=1;
   8990: out<=0;
   8991: out<=1;
   8992: out<=1;
   8993: out<=0;
   8994: out<=0;
   8995: out<=1;
   8996: out<=0;
   8997: out<=0;
   8998: out<=0;
   8999: out<=0;
   9000: out<=0;
   9001: out<=0;
   9002: out<=1;
   9003: out<=1;
   9004: out<=1;
   9005: out<=0;
   9006: out<=1;
   9007: out<=0;
   9008: out<=1;
   9009: out<=0;
   9010: out<=0;
   9011: out<=1;
   9012: out<=0;
   9013: out<=0;
   9014: out<=0;
   9015: out<=0;
   9016: out<=0;
   9017: out<=0;
   9018: out<=1;
   9019: out<=1;
   9020: out<=1;
   9021: out<=0;
   9022: out<=1;
   9023: out<=0;
   9024: out<=0;
   9025: out<=1;
   9026: out<=1;
   9027: out<=0;
   9028: out<=1;
   9029: out<=1;
   9030: out<=1;
   9031: out<=1;
   9032: out<=1;
   9033: out<=1;
   9034: out<=0;
   9035: out<=0;
   9036: out<=0;
   9037: out<=1;
   9038: out<=0;
   9039: out<=1;
   9040: out<=1;
   9041: out<=0;
   9042: out<=0;
   9043: out<=1;
   9044: out<=0;
   9045: out<=0;
   9046: out<=0;
   9047: out<=0;
   9048: out<=0;
   9049: out<=0;
   9050: out<=1;
   9051: out<=1;
   9052: out<=1;
   9053: out<=0;
   9054: out<=1;
   9055: out<=0;
   9056: out<=0;
   9057: out<=1;
   9058: out<=1;
   9059: out<=0;
   9060: out<=1;
   9061: out<=1;
   9062: out<=1;
   9063: out<=1;
   9064: out<=1;
   9065: out<=1;
   9066: out<=0;
   9067: out<=0;
   9068: out<=0;
   9069: out<=1;
   9070: out<=0;
   9071: out<=1;
   9072: out<=1;
   9073: out<=0;
   9074: out<=0;
   9075: out<=1;
   9076: out<=0;
   9077: out<=0;
   9078: out<=0;
   9079: out<=0;
   9080: out<=0;
   9081: out<=0;
   9082: out<=1;
   9083: out<=1;
   9084: out<=1;
   9085: out<=0;
   9086: out<=1;
   9087: out<=0;
   9088: out<=0;
   9089: out<=1;
   9090: out<=1;
   9091: out<=0;
   9092: out<=1;
   9093: out<=1;
   9094: out<=1;
   9095: out<=1;
   9096: out<=1;
   9097: out<=1;
   9098: out<=0;
   9099: out<=0;
   9100: out<=0;
   9101: out<=1;
   9102: out<=0;
   9103: out<=1;
   9104: out<=1;
   9105: out<=0;
   9106: out<=0;
   9107: out<=1;
   9108: out<=0;
   9109: out<=0;
   9110: out<=0;
   9111: out<=0;
   9112: out<=0;
   9113: out<=0;
   9114: out<=1;
   9115: out<=1;
   9116: out<=1;
   9117: out<=0;
   9118: out<=1;
   9119: out<=0;
   9120: out<=1;
   9121: out<=0;
   9122: out<=0;
   9123: out<=1;
   9124: out<=0;
   9125: out<=0;
   9126: out<=0;
   9127: out<=0;
   9128: out<=0;
   9129: out<=0;
   9130: out<=1;
   9131: out<=1;
   9132: out<=1;
   9133: out<=0;
   9134: out<=1;
   9135: out<=0;
   9136: out<=0;
   9137: out<=1;
   9138: out<=1;
   9139: out<=0;
   9140: out<=1;
   9141: out<=1;
   9142: out<=1;
   9143: out<=1;
   9144: out<=1;
   9145: out<=1;
   9146: out<=0;
   9147: out<=0;
   9148: out<=0;
   9149: out<=1;
   9150: out<=0;
   9151: out<=1;
   9152: out<=0;
   9153: out<=1;
   9154: out<=1;
   9155: out<=0;
   9156: out<=1;
   9157: out<=1;
   9158: out<=1;
   9159: out<=1;
   9160: out<=1;
   9161: out<=1;
   9162: out<=0;
   9163: out<=0;
   9164: out<=0;
   9165: out<=1;
   9166: out<=0;
   9167: out<=1;
   9168: out<=0;
   9169: out<=1;
   9170: out<=1;
   9171: out<=0;
   9172: out<=1;
   9173: out<=1;
   9174: out<=1;
   9175: out<=1;
   9176: out<=1;
   9177: out<=1;
   9178: out<=0;
   9179: out<=0;
   9180: out<=0;
   9181: out<=1;
   9182: out<=0;
   9183: out<=1;
   9184: out<=0;
   9185: out<=1;
   9186: out<=1;
   9187: out<=0;
   9188: out<=1;
   9189: out<=1;
   9190: out<=1;
   9191: out<=1;
   9192: out<=1;
   9193: out<=1;
   9194: out<=0;
   9195: out<=0;
   9196: out<=0;
   9197: out<=1;
   9198: out<=0;
   9199: out<=1;
   9200: out<=0;
   9201: out<=1;
   9202: out<=1;
   9203: out<=0;
   9204: out<=1;
   9205: out<=1;
   9206: out<=1;
   9207: out<=1;
   9208: out<=1;
   9209: out<=1;
   9210: out<=0;
   9211: out<=0;
   9212: out<=0;
   9213: out<=1;
   9214: out<=0;
   9215: out<=1;
   9216: out<=0;
   9217: out<=0;
   9218: out<=1;
   9219: out<=1;
   9220: out<=1;
   9221: out<=0;
   9222: out<=1;
   9223: out<=0;
   9224: out<=0;
   9225: out<=1;
   9226: out<=1;
   9227: out<=0;
   9228: out<=1;
   9229: out<=1;
   9230: out<=1;
   9231: out<=1;
   9232: out<=0;
   9233: out<=0;
   9234: out<=1;
   9235: out<=1;
   9236: out<=1;
   9237: out<=0;
   9238: out<=1;
   9239: out<=0;
   9240: out<=0;
   9241: out<=1;
   9242: out<=1;
   9243: out<=0;
   9244: out<=1;
   9245: out<=1;
   9246: out<=1;
   9247: out<=1;
   9248: out<=0;
   9249: out<=0;
   9250: out<=1;
   9251: out<=1;
   9252: out<=1;
   9253: out<=0;
   9254: out<=1;
   9255: out<=0;
   9256: out<=0;
   9257: out<=1;
   9258: out<=1;
   9259: out<=0;
   9260: out<=1;
   9261: out<=1;
   9262: out<=1;
   9263: out<=1;
   9264: out<=0;
   9265: out<=0;
   9266: out<=1;
   9267: out<=1;
   9268: out<=1;
   9269: out<=0;
   9270: out<=1;
   9271: out<=0;
   9272: out<=0;
   9273: out<=1;
   9274: out<=1;
   9275: out<=0;
   9276: out<=1;
   9277: out<=1;
   9278: out<=1;
   9279: out<=1;
   9280: out<=0;
   9281: out<=0;
   9282: out<=1;
   9283: out<=1;
   9284: out<=1;
   9285: out<=0;
   9286: out<=1;
   9287: out<=0;
   9288: out<=0;
   9289: out<=1;
   9290: out<=1;
   9291: out<=0;
   9292: out<=1;
   9293: out<=1;
   9294: out<=1;
   9295: out<=1;
   9296: out<=1;
   9297: out<=1;
   9298: out<=0;
   9299: out<=0;
   9300: out<=0;
   9301: out<=1;
   9302: out<=0;
   9303: out<=1;
   9304: out<=1;
   9305: out<=0;
   9306: out<=0;
   9307: out<=1;
   9308: out<=0;
   9309: out<=0;
   9310: out<=0;
   9311: out<=0;
   9312: out<=1;
   9313: out<=1;
   9314: out<=0;
   9315: out<=0;
   9316: out<=0;
   9317: out<=1;
   9318: out<=0;
   9319: out<=1;
   9320: out<=1;
   9321: out<=0;
   9322: out<=0;
   9323: out<=1;
   9324: out<=0;
   9325: out<=0;
   9326: out<=0;
   9327: out<=0;
   9328: out<=0;
   9329: out<=0;
   9330: out<=1;
   9331: out<=1;
   9332: out<=1;
   9333: out<=0;
   9334: out<=1;
   9335: out<=0;
   9336: out<=0;
   9337: out<=1;
   9338: out<=1;
   9339: out<=0;
   9340: out<=1;
   9341: out<=1;
   9342: out<=1;
   9343: out<=1;
   9344: out<=0;
   9345: out<=0;
   9346: out<=1;
   9347: out<=1;
   9348: out<=1;
   9349: out<=0;
   9350: out<=1;
   9351: out<=0;
   9352: out<=0;
   9353: out<=1;
   9354: out<=1;
   9355: out<=0;
   9356: out<=1;
   9357: out<=1;
   9358: out<=1;
   9359: out<=1;
   9360: out<=1;
   9361: out<=1;
   9362: out<=0;
   9363: out<=0;
   9364: out<=0;
   9365: out<=1;
   9366: out<=0;
   9367: out<=1;
   9368: out<=1;
   9369: out<=0;
   9370: out<=0;
   9371: out<=1;
   9372: out<=0;
   9373: out<=0;
   9374: out<=0;
   9375: out<=0;
   9376: out<=0;
   9377: out<=0;
   9378: out<=1;
   9379: out<=1;
   9380: out<=1;
   9381: out<=0;
   9382: out<=1;
   9383: out<=0;
   9384: out<=0;
   9385: out<=1;
   9386: out<=1;
   9387: out<=0;
   9388: out<=1;
   9389: out<=1;
   9390: out<=1;
   9391: out<=1;
   9392: out<=1;
   9393: out<=1;
   9394: out<=0;
   9395: out<=0;
   9396: out<=0;
   9397: out<=1;
   9398: out<=0;
   9399: out<=1;
   9400: out<=1;
   9401: out<=0;
   9402: out<=0;
   9403: out<=1;
   9404: out<=0;
   9405: out<=0;
   9406: out<=0;
   9407: out<=0;
   9408: out<=0;
   9409: out<=0;
   9410: out<=1;
   9411: out<=1;
   9412: out<=1;
   9413: out<=0;
   9414: out<=1;
   9415: out<=0;
   9416: out<=0;
   9417: out<=1;
   9418: out<=1;
   9419: out<=0;
   9420: out<=1;
   9421: out<=1;
   9422: out<=1;
   9423: out<=1;
   9424: out<=0;
   9425: out<=0;
   9426: out<=1;
   9427: out<=1;
   9428: out<=1;
   9429: out<=0;
   9430: out<=1;
   9431: out<=0;
   9432: out<=0;
   9433: out<=1;
   9434: out<=1;
   9435: out<=0;
   9436: out<=1;
   9437: out<=1;
   9438: out<=1;
   9439: out<=1;
   9440: out<=1;
   9441: out<=1;
   9442: out<=0;
   9443: out<=0;
   9444: out<=0;
   9445: out<=1;
   9446: out<=0;
   9447: out<=1;
   9448: out<=1;
   9449: out<=0;
   9450: out<=0;
   9451: out<=1;
   9452: out<=0;
   9453: out<=0;
   9454: out<=0;
   9455: out<=0;
   9456: out<=1;
   9457: out<=1;
   9458: out<=0;
   9459: out<=0;
   9460: out<=0;
   9461: out<=1;
   9462: out<=0;
   9463: out<=1;
   9464: out<=1;
   9465: out<=0;
   9466: out<=0;
   9467: out<=1;
   9468: out<=0;
   9469: out<=0;
   9470: out<=0;
   9471: out<=0;
   9472: out<=1;
   9473: out<=0;
   9474: out<=1;
   9475: out<=0;
   9476: out<=1;
   9477: out<=1;
   9478: out<=0;
   9479: out<=0;
   9480: out<=0;
   9481: out<=0;
   9482: out<=0;
   9483: out<=0;
   9484: out<=0;
   9485: out<=1;
   9486: out<=1;
   9487: out<=0;
   9488: out<=0;
   9489: out<=1;
   9490: out<=0;
   9491: out<=1;
   9492: out<=0;
   9493: out<=0;
   9494: out<=1;
   9495: out<=1;
   9496: out<=1;
   9497: out<=1;
   9498: out<=1;
   9499: out<=1;
   9500: out<=1;
   9501: out<=0;
   9502: out<=0;
   9503: out<=1;
   9504: out<=0;
   9505: out<=1;
   9506: out<=0;
   9507: out<=1;
   9508: out<=0;
   9509: out<=0;
   9510: out<=1;
   9511: out<=1;
   9512: out<=1;
   9513: out<=1;
   9514: out<=1;
   9515: out<=1;
   9516: out<=1;
   9517: out<=0;
   9518: out<=0;
   9519: out<=1;
   9520: out<=1;
   9521: out<=0;
   9522: out<=1;
   9523: out<=0;
   9524: out<=1;
   9525: out<=1;
   9526: out<=0;
   9527: out<=0;
   9528: out<=0;
   9529: out<=0;
   9530: out<=0;
   9531: out<=0;
   9532: out<=0;
   9533: out<=1;
   9534: out<=1;
   9535: out<=0;
   9536: out<=1;
   9537: out<=0;
   9538: out<=1;
   9539: out<=0;
   9540: out<=1;
   9541: out<=1;
   9542: out<=0;
   9543: out<=0;
   9544: out<=0;
   9545: out<=0;
   9546: out<=0;
   9547: out<=0;
   9548: out<=0;
   9549: out<=1;
   9550: out<=1;
   9551: out<=0;
   9552: out<=1;
   9553: out<=0;
   9554: out<=1;
   9555: out<=0;
   9556: out<=1;
   9557: out<=1;
   9558: out<=0;
   9559: out<=0;
   9560: out<=0;
   9561: out<=0;
   9562: out<=0;
   9563: out<=0;
   9564: out<=0;
   9565: out<=1;
   9566: out<=1;
   9567: out<=0;
   9568: out<=1;
   9569: out<=0;
   9570: out<=1;
   9571: out<=0;
   9572: out<=1;
   9573: out<=1;
   9574: out<=0;
   9575: out<=0;
   9576: out<=0;
   9577: out<=0;
   9578: out<=0;
   9579: out<=0;
   9580: out<=0;
   9581: out<=1;
   9582: out<=1;
   9583: out<=0;
   9584: out<=1;
   9585: out<=0;
   9586: out<=1;
   9587: out<=0;
   9588: out<=1;
   9589: out<=1;
   9590: out<=0;
   9591: out<=0;
   9592: out<=0;
   9593: out<=0;
   9594: out<=0;
   9595: out<=0;
   9596: out<=0;
   9597: out<=1;
   9598: out<=1;
   9599: out<=0;
   9600: out<=1;
   9601: out<=0;
   9602: out<=1;
   9603: out<=0;
   9604: out<=1;
   9605: out<=1;
   9606: out<=0;
   9607: out<=0;
   9608: out<=0;
   9609: out<=0;
   9610: out<=0;
   9611: out<=0;
   9612: out<=0;
   9613: out<=1;
   9614: out<=1;
   9615: out<=0;
   9616: out<=1;
   9617: out<=0;
   9618: out<=1;
   9619: out<=0;
   9620: out<=1;
   9621: out<=1;
   9622: out<=0;
   9623: out<=0;
   9624: out<=0;
   9625: out<=0;
   9626: out<=0;
   9627: out<=0;
   9628: out<=0;
   9629: out<=1;
   9630: out<=1;
   9631: out<=0;
   9632: out<=0;
   9633: out<=1;
   9634: out<=0;
   9635: out<=1;
   9636: out<=0;
   9637: out<=0;
   9638: out<=1;
   9639: out<=1;
   9640: out<=1;
   9641: out<=1;
   9642: out<=1;
   9643: out<=1;
   9644: out<=1;
   9645: out<=0;
   9646: out<=0;
   9647: out<=1;
   9648: out<=0;
   9649: out<=1;
   9650: out<=0;
   9651: out<=1;
   9652: out<=0;
   9653: out<=0;
   9654: out<=1;
   9655: out<=1;
   9656: out<=1;
   9657: out<=1;
   9658: out<=1;
   9659: out<=1;
   9660: out<=1;
   9661: out<=0;
   9662: out<=0;
   9663: out<=1;
   9664: out<=1;
   9665: out<=0;
   9666: out<=1;
   9667: out<=0;
   9668: out<=1;
   9669: out<=1;
   9670: out<=0;
   9671: out<=0;
   9672: out<=0;
   9673: out<=0;
   9674: out<=0;
   9675: out<=0;
   9676: out<=0;
   9677: out<=1;
   9678: out<=1;
   9679: out<=0;
   9680: out<=0;
   9681: out<=1;
   9682: out<=0;
   9683: out<=1;
   9684: out<=0;
   9685: out<=0;
   9686: out<=1;
   9687: out<=1;
   9688: out<=1;
   9689: out<=1;
   9690: out<=1;
   9691: out<=1;
   9692: out<=1;
   9693: out<=0;
   9694: out<=0;
   9695: out<=1;
   9696: out<=1;
   9697: out<=0;
   9698: out<=1;
   9699: out<=0;
   9700: out<=1;
   9701: out<=1;
   9702: out<=0;
   9703: out<=0;
   9704: out<=0;
   9705: out<=0;
   9706: out<=0;
   9707: out<=0;
   9708: out<=0;
   9709: out<=1;
   9710: out<=1;
   9711: out<=0;
   9712: out<=0;
   9713: out<=1;
   9714: out<=0;
   9715: out<=1;
   9716: out<=0;
   9717: out<=0;
   9718: out<=1;
   9719: out<=1;
   9720: out<=1;
   9721: out<=1;
   9722: out<=1;
   9723: out<=1;
   9724: out<=1;
   9725: out<=0;
   9726: out<=0;
   9727: out<=1;
   9728: out<=1;
   9729: out<=0;
   9730: out<=0;
   9731: out<=1;
   9732: out<=1;
   9733: out<=1;
   9734: out<=1;
   9735: out<=1;
   9736: out<=1;
   9737: out<=1;
   9738: out<=0;
   9739: out<=0;
   9740: out<=1;
   9741: out<=0;
   9742: out<=1;
   9743: out<=0;
   9744: out<=0;
   9745: out<=1;
   9746: out<=1;
   9747: out<=0;
   9748: out<=0;
   9749: out<=0;
   9750: out<=0;
   9751: out<=0;
   9752: out<=0;
   9753: out<=0;
   9754: out<=1;
   9755: out<=1;
   9756: out<=0;
   9757: out<=1;
   9758: out<=0;
   9759: out<=1;
   9760: out<=1;
   9761: out<=0;
   9762: out<=0;
   9763: out<=1;
   9764: out<=1;
   9765: out<=1;
   9766: out<=1;
   9767: out<=1;
   9768: out<=1;
   9769: out<=1;
   9770: out<=0;
   9771: out<=0;
   9772: out<=1;
   9773: out<=0;
   9774: out<=1;
   9775: out<=0;
   9776: out<=0;
   9777: out<=1;
   9778: out<=1;
   9779: out<=0;
   9780: out<=0;
   9781: out<=0;
   9782: out<=0;
   9783: out<=0;
   9784: out<=0;
   9785: out<=0;
   9786: out<=1;
   9787: out<=1;
   9788: out<=0;
   9789: out<=1;
   9790: out<=0;
   9791: out<=1;
   9792: out<=1;
   9793: out<=0;
   9794: out<=0;
   9795: out<=1;
   9796: out<=1;
   9797: out<=1;
   9798: out<=1;
   9799: out<=1;
   9800: out<=1;
   9801: out<=1;
   9802: out<=0;
   9803: out<=0;
   9804: out<=1;
   9805: out<=0;
   9806: out<=1;
   9807: out<=0;
   9808: out<=1;
   9809: out<=0;
   9810: out<=0;
   9811: out<=1;
   9812: out<=1;
   9813: out<=1;
   9814: out<=1;
   9815: out<=1;
   9816: out<=1;
   9817: out<=1;
   9818: out<=0;
   9819: out<=0;
   9820: out<=1;
   9821: out<=0;
   9822: out<=1;
   9823: out<=0;
   9824: out<=0;
   9825: out<=1;
   9826: out<=1;
   9827: out<=0;
   9828: out<=0;
   9829: out<=0;
   9830: out<=0;
   9831: out<=0;
   9832: out<=0;
   9833: out<=0;
   9834: out<=1;
   9835: out<=1;
   9836: out<=0;
   9837: out<=1;
   9838: out<=0;
   9839: out<=1;
   9840: out<=0;
   9841: out<=1;
   9842: out<=1;
   9843: out<=0;
   9844: out<=0;
   9845: out<=0;
   9846: out<=0;
   9847: out<=0;
   9848: out<=0;
   9849: out<=0;
   9850: out<=1;
   9851: out<=1;
   9852: out<=0;
   9853: out<=1;
   9854: out<=0;
   9855: out<=1;
   9856: out<=1;
   9857: out<=0;
   9858: out<=0;
   9859: out<=1;
   9860: out<=1;
   9861: out<=1;
   9862: out<=1;
   9863: out<=1;
   9864: out<=1;
   9865: out<=1;
   9866: out<=0;
   9867: out<=0;
   9868: out<=1;
   9869: out<=0;
   9870: out<=1;
   9871: out<=0;
   9872: out<=1;
   9873: out<=0;
   9874: out<=0;
   9875: out<=1;
   9876: out<=1;
   9877: out<=1;
   9878: out<=1;
   9879: out<=1;
   9880: out<=1;
   9881: out<=1;
   9882: out<=0;
   9883: out<=0;
   9884: out<=1;
   9885: out<=0;
   9886: out<=1;
   9887: out<=0;
   9888: out<=1;
   9889: out<=0;
   9890: out<=0;
   9891: out<=1;
   9892: out<=1;
   9893: out<=1;
   9894: out<=1;
   9895: out<=1;
   9896: out<=1;
   9897: out<=1;
   9898: out<=0;
   9899: out<=0;
   9900: out<=1;
   9901: out<=0;
   9902: out<=1;
   9903: out<=0;
   9904: out<=1;
   9905: out<=0;
   9906: out<=0;
   9907: out<=1;
   9908: out<=1;
   9909: out<=1;
   9910: out<=1;
   9911: out<=1;
   9912: out<=1;
   9913: out<=1;
   9914: out<=0;
   9915: out<=0;
   9916: out<=1;
   9917: out<=0;
   9918: out<=1;
   9919: out<=0;
   9920: out<=1;
   9921: out<=0;
   9922: out<=0;
   9923: out<=1;
   9924: out<=1;
   9925: out<=1;
   9926: out<=1;
   9927: out<=1;
   9928: out<=1;
   9929: out<=1;
   9930: out<=0;
   9931: out<=0;
   9932: out<=1;
   9933: out<=0;
   9934: out<=1;
   9935: out<=0;
   9936: out<=0;
   9937: out<=1;
   9938: out<=1;
   9939: out<=0;
   9940: out<=0;
   9941: out<=0;
   9942: out<=0;
   9943: out<=0;
   9944: out<=0;
   9945: out<=0;
   9946: out<=1;
   9947: out<=1;
   9948: out<=0;
   9949: out<=1;
   9950: out<=0;
   9951: out<=1;
   9952: out<=0;
   9953: out<=1;
   9954: out<=1;
   9955: out<=0;
   9956: out<=0;
   9957: out<=0;
   9958: out<=0;
   9959: out<=0;
   9960: out<=0;
   9961: out<=0;
   9962: out<=1;
   9963: out<=1;
   9964: out<=0;
   9965: out<=1;
   9966: out<=0;
   9967: out<=1;
   9968: out<=1;
   9969: out<=0;
   9970: out<=0;
   9971: out<=1;
   9972: out<=1;
   9973: out<=1;
   9974: out<=1;
   9975: out<=1;
   9976: out<=1;
   9977: out<=1;
   9978: out<=0;
   9979: out<=0;
   9980: out<=1;
   9981: out<=0;
   9982: out<=1;
   9983: out<=0;
   9984: out<=0;
   9985: out<=0;
   9986: out<=0;
   9987: out<=0;
   9988: out<=1;
   9989: out<=0;
   9990: out<=0;
   9991: out<=1;
   9992: out<=1;
   9993: out<=0;
   9994: out<=1;
   9995: out<=0;
   9996: out<=0;
   9997: out<=0;
   9998: out<=1;
   9999: out<=1;
   10000: out<=0;
   10001: out<=0;
   10002: out<=0;
   10003: out<=0;
   10004: out<=1;
   10005: out<=0;
   10006: out<=0;
   10007: out<=1;
   10008: out<=1;
   10009: out<=0;
   10010: out<=1;
   10011: out<=0;
   10012: out<=0;
   10013: out<=0;
   10014: out<=1;
   10015: out<=1;
   10016: out<=1;
   10017: out<=1;
   10018: out<=1;
   10019: out<=1;
   10020: out<=0;
   10021: out<=1;
   10022: out<=1;
   10023: out<=0;
   10024: out<=0;
   10025: out<=1;
   10026: out<=0;
   10027: out<=1;
   10028: out<=1;
   10029: out<=1;
   10030: out<=0;
   10031: out<=0;
   10032: out<=1;
   10033: out<=1;
   10034: out<=1;
   10035: out<=1;
   10036: out<=0;
   10037: out<=1;
   10038: out<=1;
   10039: out<=0;
   10040: out<=0;
   10041: out<=1;
   10042: out<=0;
   10043: out<=1;
   10044: out<=1;
   10045: out<=1;
   10046: out<=0;
   10047: out<=0;
   10048: out<=0;
   10049: out<=0;
   10050: out<=0;
   10051: out<=0;
   10052: out<=1;
   10053: out<=0;
   10054: out<=0;
   10055: out<=1;
   10056: out<=1;
   10057: out<=0;
   10058: out<=1;
   10059: out<=0;
   10060: out<=0;
   10061: out<=0;
   10062: out<=1;
   10063: out<=1;
   10064: out<=1;
   10065: out<=1;
   10066: out<=1;
   10067: out<=1;
   10068: out<=0;
   10069: out<=1;
   10070: out<=1;
   10071: out<=0;
   10072: out<=0;
   10073: out<=1;
   10074: out<=0;
   10075: out<=1;
   10076: out<=1;
   10077: out<=1;
   10078: out<=0;
   10079: out<=0;
   10080: out<=0;
   10081: out<=0;
   10082: out<=0;
   10083: out<=0;
   10084: out<=1;
   10085: out<=0;
   10086: out<=0;
   10087: out<=1;
   10088: out<=1;
   10089: out<=0;
   10090: out<=1;
   10091: out<=0;
   10092: out<=0;
   10093: out<=0;
   10094: out<=1;
   10095: out<=1;
   10096: out<=1;
   10097: out<=1;
   10098: out<=1;
   10099: out<=1;
   10100: out<=0;
   10101: out<=1;
   10102: out<=1;
   10103: out<=0;
   10104: out<=0;
   10105: out<=1;
   10106: out<=0;
   10107: out<=1;
   10108: out<=1;
   10109: out<=1;
   10110: out<=0;
   10111: out<=0;
   10112: out<=0;
   10113: out<=0;
   10114: out<=0;
   10115: out<=0;
   10116: out<=1;
   10117: out<=0;
   10118: out<=0;
   10119: out<=1;
   10120: out<=1;
   10121: out<=0;
   10122: out<=1;
   10123: out<=0;
   10124: out<=0;
   10125: out<=0;
   10126: out<=1;
   10127: out<=1;
   10128: out<=1;
   10129: out<=1;
   10130: out<=1;
   10131: out<=1;
   10132: out<=0;
   10133: out<=1;
   10134: out<=1;
   10135: out<=0;
   10136: out<=0;
   10137: out<=1;
   10138: out<=0;
   10139: out<=1;
   10140: out<=1;
   10141: out<=1;
   10142: out<=0;
   10143: out<=0;
   10144: out<=1;
   10145: out<=1;
   10146: out<=1;
   10147: out<=1;
   10148: out<=0;
   10149: out<=1;
   10150: out<=1;
   10151: out<=0;
   10152: out<=0;
   10153: out<=1;
   10154: out<=0;
   10155: out<=1;
   10156: out<=1;
   10157: out<=1;
   10158: out<=0;
   10159: out<=0;
   10160: out<=0;
   10161: out<=0;
   10162: out<=0;
   10163: out<=0;
   10164: out<=1;
   10165: out<=0;
   10166: out<=0;
   10167: out<=1;
   10168: out<=1;
   10169: out<=0;
   10170: out<=1;
   10171: out<=0;
   10172: out<=0;
   10173: out<=0;
   10174: out<=1;
   10175: out<=1;
   10176: out<=0;
   10177: out<=0;
   10178: out<=0;
   10179: out<=0;
   10180: out<=1;
   10181: out<=0;
   10182: out<=0;
   10183: out<=1;
   10184: out<=1;
   10185: out<=0;
   10186: out<=1;
   10187: out<=0;
   10188: out<=0;
   10189: out<=0;
   10190: out<=1;
   10191: out<=1;
   10192: out<=0;
   10193: out<=0;
   10194: out<=0;
   10195: out<=0;
   10196: out<=1;
   10197: out<=0;
   10198: out<=0;
   10199: out<=1;
   10200: out<=1;
   10201: out<=0;
   10202: out<=1;
   10203: out<=0;
   10204: out<=0;
   10205: out<=0;
   10206: out<=1;
   10207: out<=1;
   10208: out<=0;
   10209: out<=0;
   10210: out<=0;
   10211: out<=0;
   10212: out<=1;
   10213: out<=0;
   10214: out<=0;
   10215: out<=1;
   10216: out<=1;
   10217: out<=0;
   10218: out<=1;
   10219: out<=0;
   10220: out<=0;
   10221: out<=0;
   10222: out<=1;
   10223: out<=1;
   10224: out<=0;
   10225: out<=0;
   10226: out<=0;
   10227: out<=0;
   10228: out<=1;
   10229: out<=0;
   10230: out<=0;
   10231: out<=1;
   10232: out<=1;
   10233: out<=0;
   10234: out<=1;
   10235: out<=0;
   10236: out<=0;
   10237: out<=0;
   10238: out<=1;
   10239: out<=1;
   10240: out<=0;
   10241: out<=0;
   10242: out<=0;
   10243: out<=0;
   10244: out<=1;
   10245: out<=0;
   10246: out<=0;
   10247: out<=1;
   10248: out<=0;
   10249: out<=1;
   10250: out<=0;
   10251: out<=1;
   10252: out<=1;
   10253: out<=1;
   10254: out<=0;
   10255: out<=0;
   10256: out<=0;
   10257: out<=0;
   10258: out<=0;
   10259: out<=0;
   10260: out<=1;
   10261: out<=0;
   10262: out<=0;
   10263: out<=1;
   10264: out<=0;
   10265: out<=1;
   10266: out<=0;
   10267: out<=1;
   10268: out<=1;
   10269: out<=1;
   10270: out<=0;
   10271: out<=0;
   10272: out<=0;
   10273: out<=0;
   10274: out<=0;
   10275: out<=0;
   10276: out<=1;
   10277: out<=0;
   10278: out<=0;
   10279: out<=1;
   10280: out<=0;
   10281: out<=1;
   10282: out<=0;
   10283: out<=1;
   10284: out<=1;
   10285: out<=1;
   10286: out<=0;
   10287: out<=0;
   10288: out<=0;
   10289: out<=0;
   10290: out<=0;
   10291: out<=0;
   10292: out<=1;
   10293: out<=0;
   10294: out<=0;
   10295: out<=1;
   10296: out<=0;
   10297: out<=1;
   10298: out<=0;
   10299: out<=1;
   10300: out<=1;
   10301: out<=1;
   10302: out<=0;
   10303: out<=0;
   10304: out<=0;
   10305: out<=0;
   10306: out<=0;
   10307: out<=0;
   10308: out<=1;
   10309: out<=0;
   10310: out<=0;
   10311: out<=1;
   10312: out<=0;
   10313: out<=1;
   10314: out<=0;
   10315: out<=1;
   10316: out<=1;
   10317: out<=1;
   10318: out<=0;
   10319: out<=0;
   10320: out<=1;
   10321: out<=1;
   10322: out<=1;
   10323: out<=1;
   10324: out<=0;
   10325: out<=1;
   10326: out<=1;
   10327: out<=0;
   10328: out<=1;
   10329: out<=0;
   10330: out<=1;
   10331: out<=0;
   10332: out<=0;
   10333: out<=0;
   10334: out<=1;
   10335: out<=1;
   10336: out<=1;
   10337: out<=1;
   10338: out<=1;
   10339: out<=1;
   10340: out<=0;
   10341: out<=1;
   10342: out<=1;
   10343: out<=0;
   10344: out<=1;
   10345: out<=0;
   10346: out<=1;
   10347: out<=0;
   10348: out<=0;
   10349: out<=0;
   10350: out<=1;
   10351: out<=1;
   10352: out<=0;
   10353: out<=0;
   10354: out<=0;
   10355: out<=0;
   10356: out<=1;
   10357: out<=0;
   10358: out<=0;
   10359: out<=1;
   10360: out<=0;
   10361: out<=1;
   10362: out<=0;
   10363: out<=1;
   10364: out<=1;
   10365: out<=1;
   10366: out<=0;
   10367: out<=0;
   10368: out<=0;
   10369: out<=0;
   10370: out<=0;
   10371: out<=0;
   10372: out<=1;
   10373: out<=0;
   10374: out<=0;
   10375: out<=1;
   10376: out<=0;
   10377: out<=1;
   10378: out<=0;
   10379: out<=1;
   10380: out<=1;
   10381: out<=1;
   10382: out<=0;
   10383: out<=0;
   10384: out<=1;
   10385: out<=1;
   10386: out<=1;
   10387: out<=1;
   10388: out<=0;
   10389: out<=1;
   10390: out<=1;
   10391: out<=0;
   10392: out<=1;
   10393: out<=0;
   10394: out<=1;
   10395: out<=0;
   10396: out<=0;
   10397: out<=0;
   10398: out<=1;
   10399: out<=1;
   10400: out<=0;
   10401: out<=0;
   10402: out<=0;
   10403: out<=0;
   10404: out<=1;
   10405: out<=0;
   10406: out<=0;
   10407: out<=1;
   10408: out<=0;
   10409: out<=1;
   10410: out<=0;
   10411: out<=1;
   10412: out<=1;
   10413: out<=1;
   10414: out<=0;
   10415: out<=0;
   10416: out<=1;
   10417: out<=1;
   10418: out<=1;
   10419: out<=1;
   10420: out<=0;
   10421: out<=1;
   10422: out<=1;
   10423: out<=0;
   10424: out<=1;
   10425: out<=0;
   10426: out<=1;
   10427: out<=0;
   10428: out<=0;
   10429: out<=0;
   10430: out<=1;
   10431: out<=1;
   10432: out<=0;
   10433: out<=0;
   10434: out<=0;
   10435: out<=0;
   10436: out<=1;
   10437: out<=0;
   10438: out<=0;
   10439: out<=1;
   10440: out<=0;
   10441: out<=1;
   10442: out<=0;
   10443: out<=1;
   10444: out<=1;
   10445: out<=1;
   10446: out<=0;
   10447: out<=0;
   10448: out<=0;
   10449: out<=0;
   10450: out<=0;
   10451: out<=0;
   10452: out<=1;
   10453: out<=0;
   10454: out<=0;
   10455: out<=1;
   10456: out<=0;
   10457: out<=1;
   10458: out<=0;
   10459: out<=1;
   10460: out<=1;
   10461: out<=1;
   10462: out<=0;
   10463: out<=0;
   10464: out<=1;
   10465: out<=1;
   10466: out<=1;
   10467: out<=1;
   10468: out<=0;
   10469: out<=1;
   10470: out<=1;
   10471: out<=0;
   10472: out<=1;
   10473: out<=0;
   10474: out<=1;
   10475: out<=0;
   10476: out<=0;
   10477: out<=0;
   10478: out<=1;
   10479: out<=1;
   10480: out<=1;
   10481: out<=1;
   10482: out<=1;
   10483: out<=1;
   10484: out<=0;
   10485: out<=1;
   10486: out<=1;
   10487: out<=0;
   10488: out<=1;
   10489: out<=0;
   10490: out<=1;
   10491: out<=0;
   10492: out<=0;
   10493: out<=0;
   10494: out<=1;
   10495: out<=1;
   10496: out<=1;
   10497: out<=0;
   10498: out<=0;
   10499: out<=1;
   10500: out<=1;
   10501: out<=1;
   10502: out<=1;
   10503: out<=1;
   10504: out<=0;
   10505: out<=0;
   10506: out<=1;
   10507: out<=1;
   10508: out<=0;
   10509: out<=1;
   10510: out<=0;
   10511: out<=1;
   10512: out<=0;
   10513: out<=1;
   10514: out<=1;
   10515: out<=0;
   10516: out<=0;
   10517: out<=0;
   10518: out<=0;
   10519: out<=0;
   10520: out<=1;
   10521: out<=1;
   10522: out<=0;
   10523: out<=0;
   10524: out<=1;
   10525: out<=0;
   10526: out<=1;
   10527: out<=0;
   10528: out<=0;
   10529: out<=1;
   10530: out<=1;
   10531: out<=0;
   10532: out<=0;
   10533: out<=0;
   10534: out<=0;
   10535: out<=0;
   10536: out<=1;
   10537: out<=1;
   10538: out<=0;
   10539: out<=0;
   10540: out<=1;
   10541: out<=0;
   10542: out<=1;
   10543: out<=0;
   10544: out<=1;
   10545: out<=0;
   10546: out<=0;
   10547: out<=1;
   10548: out<=1;
   10549: out<=1;
   10550: out<=1;
   10551: out<=1;
   10552: out<=0;
   10553: out<=0;
   10554: out<=1;
   10555: out<=1;
   10556: out<=0;
   10557: out<=1;
   10558: out<=0;
   10559: out<=1;
   10560: out<=1;
   10561: out<=0;
   10562: out<=0;
   10563: out<=1;
   10564: out<=1;
   10565: out<=1;
   10566: out<=1;
   10567: out<=1;
   10568: out<=0;
   10569: out<=0;
   10570: out<=1;
   10571: out<=1;
   10572: out<=0;
   10573: out<=1;
   10574: out<=0;
   10575: out<=1;
   10576: out<=1;
   10577: out<=0;
   10578: out<=0;
   10579: out<=1;
   10580: out<=1;
   10581: out<=1;
   10582: out<=1;
   10583: out<=1;
   10584: out<=0;
   10585: out<=0;
   10586: out<=1;
   10587: out<=1;
   10588: out<=0;
   10589: out<=1;
   10590: out<=0;
   10591: out<=1;
   10592: out<=1;
   10593: out<=0;
   10594: out<=0;
   10595: out<=1;
   10596: out<=1;
   10597: out<=1;
   10598: out<=1;
   10599: out<=1;
   10600: out<=0;
   10601: out<=0;
   10602: out<=1;
   10603: out<=1;
   10604: out<=0;
   10605: out<=1;
   10606: out<=0;
   10607: out<=1;
   10608: out<=1;
   10609: out<=0;
   10610: out<=0;
   10611: out<=1;
   10612: out<=1;
   10613: out<=1;
   10614: out<=1;
   10615: out<=1;
   10616: out<=0;
   10617: out<=0;
   10618: out<=1;
   10619: out<=1;
   10620: out<=0;
   10621: out<=1;
   10622: out<=0;
   10623: out<=1;
   10624: out<=1;
   10625: out<=0;
   10626: out<=0;
   10627: out<=1;
   10628: out<=1;
   10629: out<=1;
   10630: out<=1;
   10631: out<=1;
   10632: out<=0;
   10633: out<=0;
   10634: out<=1;
   10635: out<=1;
   10636: out<=0;
   10637: out<=1;
   10638: out<=0;
   10639: out<=1;
   10640: out<=1;
   10641: out<=0;
   10642: out<=0;
   10643: out<=1;
   10644: out<=1;
   10645: out<=1;
   10646: out<=1;
   10647: out<=1;
   10648: out<=0;
   10649: out<=0;
   10650: out<=1;
   10651: out<=1;
   10652: out<=0;
   10653: out<=1;
   10654: out<=0;
   10655: out<=1;
   10656: out<=0;
   10657: out<=1;
   10658: out<=1;
   10659: out<=0;
   10660: out<=0;
   10661: out<=0;
   10662: out<=0;
   10663: out<=0;
   10664: out<=1;
   10665: out<=1;
   10666: out<=0;
   10667: out<=0;
   10668: out<=1;
   10669: out<=0;
   10670: out<=1;
   10671: out<=0;
   10672: out<=0;
   10673: out<=1;
   10674: out<=1;
   10675: out<=0;
   10676: out<=0;
   10677: out<=0;
   10678: out<=0;
   10679: out<=0;
   10680: out<=1;
   10681: out<=1;
   10682: out<=0;
   10683: out<=0;
   10684: out<=1;
   10685: out<=0;
   10686: out<=1;
   10687: out<=0;
   10688: out<=1;
   10689: out<=0;
   10690: out<=0;
   10691: out<=1;
   10692: out<=1;
   10693: out<=1;
   10694: out<=1;
   10695: out<=1;
   10696: out<=0;
   10697: out<=0;
   10698: out<=1;
   10699: out<=1;
   10700: out<=0;
   10701: out<=1;
   10702: out<=0;
   10703: out<=1;
   10704: out<=0;
   10705: out<=1;
   10706: out<=1;
   10707: out<=0;
   10708: out<=0;
   10709: out<=0;
   10710: out<=0;
   10711: out<=0;
   10712: out<=1;
   10713: out<=1;
   10714: out<=0;
   10715: out<=0;
   10716: out<=1;
   10717: out<=0;
   10718: out<=1;
   10719: out<=0;
   10720: out<=1;
   10721: out<=0;
   10722: out<=0;
   10723: out<=1;
   10724: out<=1;
   10725: out<=1;
   10726: out<=1;
   10727: out<=1;
   10728: out<=0;
   10729: out<=0;
   10730: out<=1;
   10731: out<=1;
   10732: out<=0;
   10733: out<=1;
   10734: out<=0;
   10735: out<=1;
   10736: out<=0;
   10737: out<=1;
   10738: out<=1;
   10739: out<=0;
   10740: out<=0;
   10741: out<=0;
   10742: out<=0;
   10743: out<=0;
   10744: out<=1;
   10745: out<=1;
   10746: out<=0;
   10747: out<=0;
   10748: out<=1;
   10749: out<=0;
   10750: out<=1;
   10751: out<=0;
   10752: out<=0;
   10753: out<=1;
   10754: out<=0;
   10755: out<=1;
   10756: out<=0;
   10757: out<=0;
   10758: out<=1;
   10759: out<=1;
   10760: out<=0;
   10761: out<=0;
   10762: out<=0;
   10763: out<=0;
   10764: out<=0;
   10765: out<=1;
   10766: out<=1;
   10767: out<=0;
   10768: out<=1;
   10769: out<=0;
   10770: out<=1;
   10771: out<=0;
   10772: out<=1;
   10773: out<=1;
   10774: out<=0;
   10775: out<=0;
   10776: out<=1;
   10777: out<=1;
   10778: out<=1;
   10779: out<=1;
   10780: out<=1;
   10781: out<=0;
   10782: out<=0;
   10783: out<=1;
   10784: out<=0;
   10785: out<=1;
   10786: out<=0;
   10787: out<=1;
   10788: out<=0;
   10789: out<=0;
   10790: out<=1;
   10791: out<=1;
   10792: out<=0;
   10793: out<=0;
   10794: out<=0;
   10795: out<=0;
   10796: out<=0;
   10797: out<=1;
   10798: out<=1;
   10799: out<=0;
   10800: out<=1;
   10801: out<=0;
   10802: out<=1;
   10803: out<=0;
   10804: out<=1;
   10805: out<=1;
   10806: out<=0;
   10807: out<=0;
   10808: out<=1;
   10809: out<=1;
   10810: out<=1;
   10811: out<=1;
   10812: out<=1;
   10813: out<=0;
   10814: out<=0;
   10815: out<=1;
   10816: out<=0;
   10817: out<=1;
   10818: out<=0;
   10819: out<=1;
   10820: out<=0;
   10821: out<=0;
   10822: out<=1;
   10823: out<=1;
   10824: out<=0;
   10825: out<=0;
   10826: out<=0;
   10827: out<=0;
   10828: out<=0;
   10829: out<=1;
   10830: out<=1;
   10831: out<=0;
   10832: out<=0;
   10833: out<=1;
   10834: out<=0;
   10835: out<=1;
   10836: out<=0;
   10837: out<=0;
   10838: out<=1;
   10839: out<=1;
   10840: out<=0;
   10841: out<=0;
   10842: out<=0;
   10843: out<=0;
   10844: out<=0;
   10845: out<=1;
   10846: out<=1;
   10847: out<=0;
   10848: out<=1;
   10849: out<=0;
   10850: out<=1;
   10851: out<=0;
   10852: out<=1;
   10853: out<=1;
   10854: out<=0;
   10855: out<=0;
   10856: out<=1;
   10857: out<=1;
   10858: out<=1;
   10859: out<=1;
   10860: out<=1;
   10861: out<=0;
   10862: out<=0;
   10863: out<=1;
   10864: out<=1;
   10865: out<=0;
   10866: out<=1;
   10867: out<=0;
   10868: out<=1;
   10869: out<=1;
   10870: out<=0;
   10871: out<=0;
   10872: out<=1;
   10873: out<=1;
   10874: out<=1;
   10875: out<=1;
   10876: out<=1;
   10877: out<=0;
   10878: out<=0;
   10879: out<=1;
   10880: out<=0;
   10881: out<=1;
   10882: out<=0;
   10883: out<=1;
   10884: out<=0;
   10885: out<=0;
   10886: out<=1;
   10887: out<=1;
   10888: out<=0;
   10889: out<=0;
   10890: out<=0;
   10891: out<=0;
   10892: out<=0;
   10893: out<=1;
   10894: out<=1;
   10895: out<=0;
   10896: out<=0;
   10897: out<=1;
   10898: out<=0;
   10899: out<=1;
   10900: out<=0;
   10901: out<=0;
   10902: out<=1;
   10903: out<=1;
   10904: out<=0;
   10905: out<=0;
   10906: out<=0;
   10907: out<=0;
   10908: out<=0;
   10909: out<=1;
   10910: out<=1;
   10911: out<=0;
   10912: out<=0;
   10913: out<=1;
   10914: out<=0;
   10915: out<=1;
   10916: out<=0;
   10917: out<=0;
   10918: out<=1;
   10919: out<=1;
   10920: out<=0;
   10921: out<=0;
   10922: out<=0;
   10923: out<=0;
   10924: out<=0;
   10925: out<=1;
   10926: out<=1;
   10927: out<=0;
   10928: out<=0;
   10929: out<=1;
   10930: out<=0;
   10931: out<=1;
   10932: out<=0;
   10933: out<=0;
   10934: out<=1;
   10935: out<=1;
   10936: out<=0;
   10937: out<=0;
   10938: out<=0;
   10939: out<=0;
   10940: out<=0;
   10941: out<=1;
   10942: out<=1;
   10943: out<=0;
   10944: out<=0;
   10945: out<=1;
   10946: out<=0;
   10947: out<=1;
   10948: out<=0;
   10949: out<=0;
   10950: out<=1;
   10951: out<=1;
   10952: out<=0;
   10953: out<=0;
   10954: out<=0;
   10955: out<=0;
   10956: out<=0;
   10957: out<=1;
   10958: out<=1;
   10959: out<=0;
   10960: out<=1;
   10961: out<=0;
   10962: out<=1;
   10963: out<=0;
   10964: out<=1;
   10965: out<=1;
   10966: out<=0;
   10967: out<=0;
   10968: out<=1;
   10969: out<=1;
   10970: out<=1;
   10971: out<=1;
   10972: out<=1;
   10973: out<=0;
   10974: out<=0;
   10975: out<=1;
   10976: out<=1;
   10977: out<=0;
   10978: out<=1;
   10979: out<=0;
   10980: out<=1;
   10981: out<=1;
   10982: out<=0;
   10983: out<=0;
   10984: out<=1;
   10985: out<=1;
   10986: out<=1;
   10987: out<=1;
   10988: out<=1;
   10989: out<=0;
   10990: out<=0;
   10991: out<=1;
   10992: out<=0;
   10993: out<=1;
   10994: out<=0;
   10995: out<=1;
   10996: out<=0;
   10997: out<=0;
   10998: out<=1;
   10999: out<=1;
   11000: out<=0;
   11001: out<=0;
   11002: out<=0;
   11003: out<=0;
   11004: out<=0;
   11005: out<=1;
   11006: out<=1;
   11007: out<=0;
   11008: out<=1;
   11009: out<=1;
   11010: out<=0;
   11011: out<=0;
   11012: out<=0;
   11013: out<=1;
   11014: out<=0;
   11015: out<=1;
   11016: out<=0;
   11017: out<=1;
   11018: out<=1;
   11019: out<=0;
   11020: out<=1;
   11021: out<=1;
   11022: out<=1;
   11023: out<=1;
   11024: out<=1;
   11025: out<=1;
   11026: out<=0;
   11027: out<=0;
   11028: out<=0;
   11029: out<=1;
   11030: out<=0;
   11031: out<=1;
   11032: out<=0;
   11033: out<=1;
   11034: out<=1;
   11035: out<=0;
   11036: out<=1;
   11037: out<=1;
   11038: out<=1;
   11039: out<=1;
   11040: out<=0;
   11041: out<=0;
   11042: out<=1;
   11043: out<=1;
   11044: out<=1;
   11045: out<=0;
   11046: out<=1;
   11047: out<=0;
   11048: out<=1;
   11049: out<=0;
   11050: out<=0;
   11051: out<=1;
   11052: out<=0;
   11053: out<=0;
   11054: out<=0;
   11055: out<=0;
   11056: out<=0;
   11057: out<=0;
   11058: out<=1;
   11059: out<=1;
   11060: out<=1;
   11061: out<=0;
   11062: out<=1;
   11063: out<=0;
   11064: out<=1;
   11065: out<=0;
   11066: out<=0;
   11067: out<=1;
   11068: out<=0;
   11069: out<=0;
   11070: out<=0;
   11071: out<=0;
   11072: out<=1;
   11073: out<=1;
   11074: out<=0;
   11075: out<=0;
   11076: out<=0;
   11077: out<=1;
   11078: out<=0;
   11079: out<=1;
   11080: out<=0;
   11081: out<=1;
   11082: out<=1;
   11083: out<=0;
   11084: out<=1;
   11085: out<=1;
   11086: out<=1;
   11087: out<=1;
   11088: out<=0;
   11089: out<=0;
   11090: out<=1;
   11091: out<=1;
   11092: out<=1;
   11093: out<=0;
   11094: out<=1;
   11095: out<=0;
   11096: out<=1;
   11097: out<=0;
   11098: out<=0;
   11099: out<=1;
   11100: out<=0;
   11101: out<=0;
   11102: out<=0;
   11103: out<=0;
   11104: out<=1;
   11105: out<=1;
   11106: out<=0;
   11107: out<=0;
   11108: out<=0;
   11109: out<=1;
   11110: out<=0;
   11111: out<=1;
   11112: out<=0;
   11113: out<=1;
   11114: out<=1;
   11115: out<=0;
   11116: out<=1;
   11117: out<=1;
   11118: out<=1;
   11119: out<=1;
   11120: out<=0;
   11121: out<=0;
   11122: out<=1;
   11123: out<=1;
   11124: out<=1;
   11125: out<=0;
   11126: out<=1;
   11127: out<=0;
   11128: out<=1;
   11129: out<=0;
   11130: out<=0;
   11131: out<=1;
   11132: out<=0;
   11133: out<=0;
   11134: out<=0;
   11135: out<=0;
   11136: out<=1;
   11137: out<=1;
   11138: out<=0;
   11139: out<=0;
   11140: out<=0;
   11141: out<=1;
   11142: out<=0;
   11143: out<=1;
   11144: out<=0;
   11145: out<=1;
   11146: out<=1;
   11147: out<=0;
   11148: out<=1;
   11149: out<=1;
   11150: out<=1;
   11151: out<=1;
   11152: out<=0;
   11153: out<=0;
   11154: out<=1;
   11155: out<=1;
   11156: out<=1;
   11157: out<=0;
   11158: out<=1;
   11159: out<=0;
   11160: out<=1;
   11161: out<=0;
   11162: out<=0;
   11163: out<=1;
   11164: out<=0;
   11165: out<=0;
   11166: out<=0;
   11167: out<=0;
   11168: out<=0;
   11169: out<=0;
   11170: out<=1;
   11171: out<=1;
   11172: out<=1;
   11173: out<=0;
   11174: out<=1;
   11175: out<=0;
   11176: out<=1;
   11177: out<=0;
   11178: out<=0;
   11179: out<=1;
   11180: out<=0;
   11181: out<=0;
   11182: out<=0;
   11183: out<=0;
   11184: out<=1;
   11185: out<=1;
   11186: out<=0;
   11187: out<=0;
   11188: out<=0;
   11189: out<=1;
   11190: out<=0;
   11191: out<=1;
   11192: out<=0;
   11193: out<=1;
   11194: out<=1;
   11195: out<=0;
   11196: out<=1;
   11197: out<=1;
   11198: out<=1;
   11199: out<=1;
   11200: out<=1;
   11201: out<=1;
   11202: out<=0;
   11203: out<=0;
   11204: out<=0;
   11205: out<=1;
   11206: out<=0;
   11207: out<=1;
   11208: out<=0;
   11209: out<=1;
   11210: out<=1;
   11211: out<=0;
   11212: out<=1;
   11213: out<=1;
   11214: out<=1;
   11215: out<=1;
   11216: out<=1;
   11217: out<=1;
   11218: out<=0;
   11219: out<=0;
   11220: out<=0;
   11221: out<=1;
   11222: out<=0;
   11223: out<=1;
   11224: out<=0;
   11225: out<=1;
   11226: out<=1;
   11227: out<=0;
   11228: out<=1;
   11229: out<=1;
   11230: out<=1;
   11231: out<=1;
   11232: out<=1;
   11233: out<=1;
   11234: out<=0;
   11235: out<=0;
   11236: out<=0;
   11237: out<=1;
   11238: out<=0;
   11239: out<=1;
   11240: out<=0;
   11241: out<=1;
   11242: out<=1;
   11243: out<=0;
   11244: out<=1;
   11245: out<=1;
   11246: out<=1;
   11247: out<=1;
   11248: out<=1;
   11249: out<=1;
   11250: out<=0;
   11251: out<=0;
   11252: out<=0;
   11253: out<=1;
   11254: out<=0;
   11255: out<=1;
   11256: out<=0;
   11257: out<=1;
   11258: out<=1;
   11259: out<=0;
   11260: out<=1;
   11261: out<=1;
   11262: out<=1;
   11263: out<=1;
   11264: out<=0;
   11265: out<=1;
   11266: out<=1;
   11267: out<=0;
   11268: out<=1;
   11269: out<=1;
   11270: out<=1;
   11271: out<=1;
   11272: out<=0;
   11273: out<=0;
   11274: out<=1;
   11275: out<=1;
   11276: out<=1;
   11277: out<=0;
   11278: out<=1;
   11279: out<=0;
   11280: out<=0;
   11281: out<=1;
   11282: out<=1;
   11283: out<=0;
   11284: out<=1;
   11285: out<=1;
   11286: out<=1;
   11287: out<=1;
   11288: out<=0;
   11289: out<=0;
   11290: out<=1;
   11291: out<=1;
   11292: out<=1;
   11293: out<=0;
   11294: out<=1;
   11295: out<=0;
   11296: out<=0;
   11297: out<=1;
   11298: out<=1;
   11299: out<=0;
   11300: out<=1;
   11301: out<=1;
   11302: out<=1;
   11303: out<=1;
   11304: out<=0;
   11305: out<=0;
   11306: out<=1;
   11307: out<=1;
   11308: out<=1;
   11309: out<=0;
   11310: out<=1;
   11311: out<=0;
   11312: out<=0;
   11313: out<=1;
   11314: out<=1;
   11315: out<=0;
   11316: out<=1;
   11317: out<=1;
   11318: out<=1;
   11319: out<=1;
   11320: out<=0;
   11321: out<=0;
   11322: out<=1;
   11323: out<=1;
   11324: out<=1;
   11325: out<=0;
   11326: out<=1;
   11327: out<=0;
   11328: out<=0;
   11329: out<=1;
   11330: out<=1;
   11331: out<=0;
   11332: out<=1;
   11333: out<=1;
   11334: out<=1;
   11335: out<=1;
   11336: out<=0;
   11337: out<=0;
   11338: out<=1;
   11339: out<=1;
   11340: out<=1;
   11341: out<=0;
   11342: out<=1;
   11343: out<=0;
   11344: out<=1;
   11345: out<=0;
   11346: out<=0;
   11347: out<=1;
   11348: out<=0;
   11349: out<=0;
   11350: out<=0;
   11351: out<=0;
   11352: out<=1;
   11353: out<=1;
   11354: out<=0;
   11355: out<=0;
   11356: out<=0;
   11357: out<=1;
   11358: out<=0;
   11359: out<=1;
   11360: out<=1;
   11361: out<=0;
   11362: out<=0;
   11363: out<=1;
   11364: out<=0;
   11365: out<=0;
   11366: out<=0;
   11367: out<=0;
   11368: out<=1;
   11369: out<=1;
   11370: out<=0;
   11371: out<=0;
   11372: out<=0;
   11373: out<=1;
   11374: out<=0;
   11375: out<=1;
   11376: out<=0;
   11377: out<=1;
   11378: out<=1;
   11379: out<=0;
   11380: out<=1;
   11381: out<=1;
   11382: out<=1;
   11383: out<=1;
   11384: out<=0;
   11385: out<=0;
   11386: out<=1;
   11387: out<=1;
   11388: out<=1;
   11389: out<=0;
   11390: out<=1;
   11391: out<=0;
   11392: out<=0;
   11393: out<=1;
   11394: out<=1;
   11395: out<=0;
   11396: out<=1;
   11397: out<=1;
   11398: out<=1;
   11399: out<=1;
   11400: out<=0;
   11401: out<=0;
   11402: out<=1;
   11403: out<=1;
   11404: out<=1;
   11405: out<=0;
   11406: out<=1;
   11407: out<=0;
   11408: out<=1;
   11409: out<=0;
   11410: out<=0;
   11411: out<=1;
   11412: out<=0;
   11413: out<=0;
   11414: out<=0;
   11415: out<=0;
   11416: out<=1;
   11417: out<=1;
   11418: out<=0;
   11419: out<=0;
   11420: out<=0;
   11421: out<=1;
   11422: out<=0;
   11423: out<=1;
   11424: out<=0;
   11425: out<=1;
   11426: out<=1;
   11427: out<=0;
   11428: out<=1;
   11429: out<=1;
   11430: out<=1;
   11431: out<=1;
   11432: out<=0;
   11433: out<=0;
   11434: out<=1;
   11435: out<=1;
   11436: out<=1;
   11437: out<=0;
   11438: out<=1;
   11439: out<=0;
   11440: out<=1;
   11441: out<=0;
   11442: out<=0;
   11443: out<=1;
   11444: out<=0;
   11445: out<=0;
   11446: out<=0;
   11447: out<=0;
   11448: out<=1;
   11449: out<=1;
   11450: out<=0;
   11451: out<=0;
   11452: out<=0;
   11453: out<=1;
   11454: out<=0;
   11455: out<=1;
   11456: out<=0;
   11457: out<=1;
   11458: out<=1;
   11459: out<=0;
   11460: out<=1;
   11461: out<=1;
   11462: out<=1;
   11463: out<=1;
   11464: out<=0;
   11465: out<=0;
   11466: out<=1;
   11467: out<=1;
   11468: out<=1;
   11469: out<=0;
   11470: out<=1;
   11471: out<=0;
   11472: out<=0;
   11473: out<=1;
   11474: out<=1;
   11475: out<=0;
   11476: out<=1;
   11477: out<=1;
   11478: out<=1;
   11479: out<=1;
   11480: out<=0;
   11481: out<=0;
   11482: out<=1;
   11483: out<=1;
   11484: out<=1;
   11485: out<=0;
   11486: out<=1;
   11487: out<=0;
   11488: out<=1;
   11489: out<=0;
   11490: out<=0;
   11491: out<=1;
   11492: out<=0;
   11493: out<=0;
   11494: out<=0;
   11495: out<=0;
   11496: out<=1;
   11497: out<=1;
   11498: out<=0;
   11499: out<=0;
   11500: out<=0;
   11501: out<=1;
   11502: out<=0;
   11503: out<=1;
   11504: out<=1;
   11505: out<=0;
   11506: out<=0;
   11507: out<=1;
   11508: out<=0;
   11509: out<=0;
   11510: out<=0;
   11511: out<=0;
   11512: out<=1;
   11513: out<=1;
   11514: out<=0;
   11515: out<=0;
   11516: out<=0;
   11517: out<=1;
   11518: out<=0;
   11519: out<=1;
   11520: out<=0;
   11521: out<=0;
   11522: out<=0;
   11523: out<=0;
   11524: out<=0;
   11525: out<=1;
   11526: out<=1;
   11527: out<=0;
   11528: out<=1;
   11529: out<=0;
   11530: out<=1;
   11531: out<=0;
   11532: out<=1;
   11533: out<=1;
   11534: out<=0;
   11535: out<=0;
   11536: out<=1;
   11537: out<=1;
   11538: out<=1;
   11539: out<=1;
   11540: out<=1;
   11541: out<=0;
   11542: out<=0;
   11543: out<=1;
   11544: out<=0;
   11545: out<=1;
   11546: out<=0;
   11547: out<=1;
   11548: out<=0;
   11549: out<=0;
   11550: out<=1;
   11551: out<=1;
   11552: out<=1;
   11553: out<=1;
   11554: out<=1;
   11555: out<=1;
   11556: out<=1;
   11557: out<=0;
   11558: out<=0;
   11559: out<=1;
   11560: out<=0;
   11561: out<=1;
   11562: out<=0;
   11563: out<=1;
   11564: out<=0;
   11565: out<=0;
   11566: out<=1;
   11567: out<=1;
   11568: out<=0;
   11569: out<=0;
   11570: out<=0;
   11571: out<=0;
   11572: out<=0;
   11573: out<=1;
   11574: out<=1;
   11575: out<=0;
   11576: out<=1;
   11577: out<=0;
   11578: out<=1;
   11579: out<=0;
   11580: out<=1;
   11581: out<=1;
   11582: out<=0;
   11583: out<=0;
   11584: out<=0;
   11585: out<=0;
   11586: out<=0;
   11587: out<=0;
   11588: out<=0;
   11589: out<=1;
   11590: out<=1;
   11591: out<=0;
   11592: out<=1;
   11593: out<=0;
   11594: out<=1;
   11595: out<=0;
   11596: out<=1;
   11597: out<=1;
   11598: out<=0;
   11599: out<=0;
   11600: out<=0;
   11601: out<=0;
   11602: out<=0;
   11603: out<=0;
   11604: out<=0;
   11605: out<=1;
   11606: out<=1;
   11607: out<=0;
   11608: out<=1;
   11609: out<=0;
   11610: out<=1;
   11611: out<=0;
   11612: out<=1;
   11613: out<=1;
   11614: out<=0;
   11615: out<=0;
   11616: out<=0;
   11617: out<=0;
   11618: out<=0;
   11619: out<=0;
   11620: out<=0;
   11621: out<=1;
   11622: out<=1;
   11623: out<=0;
   11624: out<=1;
   11625: out<=0;
   11626: out<=1;
   11627: out<=0;
   11628: out<=1;
   11629: out<=1;
   11630: out<=0;
   11631: out<=0;
   11632: out<=0;
   11633: out<=0;
   11634: out<=0;
   11635: out<=0;
   11636: out<=0;
   11637: out<=1;
   11638: out<=1;
   11639: out<=0;
   11640: out<=1;
   11641: out<=0;
   11642: out<=1;
   11643: out<=0;
   11644: out<=1;
   11645: out<=1;
   11646: out<=0;
   11647: out<=0;
   11648: out<=0;
   11649: out<=0;
   11650: out<=0;
   11651: out<=0;
   11652: out<=0;
   11653: out<=1;
   11654: out<=1;
   11655: out<=0;
   11656: out<=1;
   11657: out<=0;
   11658: out<=1;
   11659: out<=0;
   11660: out<=1;
   11661: out<=1;
   11662: out<=0;
   11663: out<=0;
   11664: out<=0;
   11665: out<=0;
   11666: out<=0;
   11667: out<=0;
   11668: out<=0;
   11669: out<=1;
   11670: out<=1;
   11671: out<=0;
   11672: out<=1;
   11673: out<=0;
   11674: out<=1;
   11675: out<=0;
   11676: out<=1;
   11677: out<=1;
   11678: out<=0;
   11679: out<=0;
   11680: out<=1;
   11681: out<=1;
   11682: out<=1;
   11683: out<=1;
   11684: out<=1;
   11685: out<=0;
   11686: out<=0;
   11687: out<=1;
   11688: out<=0;
   11689: out<=1;
   11690: out<=0;
   11691: out<=1;
   11692: out<=0;
   11693: out<=0;
   11694: out<=1;
   11695: out<=1;
   11696: out<=1;
   11697: out<=1;
   11698: out<=1;
   11699: out<=1;
   11700: out<=1;
   11701: out<=0;
   11702: out<=0;
   11703: out<=1;
   11704: out<=0;
   11705: out<=1;
   11706: out<=0;
   11707: out<=1;
   11708: out<=0;
   11709: out<=0;
   11710: out<=1;
   11711: out<=1;
   11712: out<=0;
   11713: out<=0;
   11714: out<=0;
   11715: out<=0;
   11716: out<=0;
   11717: out<=1;
   11718: out<=1;
   11719: out<=0;
   11720: out<=1;
   11721: out<=0;
   11722: out<=1;
   11723: out<=0;
   11724: out<=1;
   11725: out<=1;
   11726: out<=0;
   11727: out<=0;
   11728: out<=1;
   11729: out<=1;
   11730: out<=1;
   11731: out<=1;
   11732: out<=1;
   11733: out<=0;
   11734: out<=0;
   11735: out<=1;
   11736: out<=0;
   11737: out<=1;
   11738: out<=0;
   11739: out<=1;
   11740: out<=0;
   11741: out<=0;
   11742: out<=1;
   11743: out<=1;
   11744: out<=0;
   11745: out<=0;
   11746: out<=0;
   11747: out<=0;
   11748: out<=0;
   11749: out<=1;
   11750: out<=1;
   11751: out<=0;
   11752: out<=1;
   11753: out<=0;
   11754: out<=1;
   11755: out<=0;
   11756: out<=1;
   11757: out<=1;
   11758: out<=0;
   11759: out<=0;
   11760: out<=1;
   11761: out<=1;
   11762: out<=1;
   11763: out<=1;
   11764: out<=1;
   11765: out<=0;
   11766: out<=0;
   11767: out<=1;
   11768: out<=0;
   11769: out<=1;
   11770: out<=0;
   11771: out<=1;
   11772: out<=0;
   11773: out<=0;
   11774: out<=1;
   11775: out<=1;
   11776: out<=1;
   11777: out<=1;
   11778: out<=0;
   11779: out<=0;
   11780: out<=1;
   11781: out<=0;
   11782: out<=1;
   11783: out<=0;
   11784: out<=1;
   11785: out<=0;
   11786: out<=0;
   11787: out<=1;
   11788: out<=1;
   11789: out<=1;
   11790: out<=1;
   11791: out<=1;
   11792: out<=0;
   11793: out<=0;
   11794: out<=1;
   11795: out<=1;
   11796: out<=0;
   11797: out<=1;
   11798: out<=0;
   11799: out<=1;
   11800: out<=0;
   11801: out<=1;
   11802: out<=1;
   11803: out<=0;
   11804: out<=0;
   11805: out<=0;
   11806: out<=0;
   11807: out<=0;
   11808: out<=1;
   11809: out<=1;
   11810: out<=0;
   11811: out<=0;
   11812: out<=1;
   11813: out<=0;
   11814: out<=1;
   11815: out<=0;
   11816: out<=1;
   11817: out<=0;
   11818: out<=0;
   11819: out<=1;
   11820: out<=1;
   11821: out<=1;
   11822: out<=1;
   11823: out<=1;
   11824: out<=0;
   11825: out<=0;
   11826: out<=1;
   11827: out<=1;
   11828: out<=0;
   11829: out<=1;
   11830: out<=0;
   11831: out<=1;
   11832: out<=0;
   11833: out<=1;
   11834: out<=1;
   11835: out<=0;
   11836: out<=0;
   11837: out<=0;
   11838: out<=0;
   11839: out<=0;
   11840: out<=1;
   11841: out<=1;
   11842: out<=0;
   11843: out<=0;
   11844: out<=1;
   11845: out<=0;
   11846: out<=1;
   11847: out<=0;
   11848: out<=1;
   11849: out<=0;
   11850: out<=0;
   11851: out<=1;
   11852: out<=1;
   11853: out<=1;
   11854: out<=1;
   11855: out<=1;
   11856: out<=1;
   11857: out<=1;
   11858: out<=0;
   11859: out<=0;
   11860: out<=1;
   11861: out<=0;
   11862: out<=1;
   11863: out<=0;
   11864: out<=1;
   11865: out<=0;
   11866: out<=0;
   11867: out<=1;
   11868: out<=1;
   11869: out<=1;
   11870: out<=1;
   11871: out<=1;
   11872: out<=0;
   11873: out<=0;
   11874: out<=1;
   11875: out<=1;
   11876: out<=0;
   11877: out<=1;
   11878: out<=0;
   11879: out<=1;
   11880: out<=0;
   11881: out<=1;
   11882: out<=1;
   11883: out<=0;
   11884: out<=0;
   11885: out<=0;
   11886: out<=0;
   11887: out<=0;
   11888: out<=0;
   11889: out<=0;
   11890: out<=1;
   11891: out<=1;
   11892: out<=0;
   11893: out<=1;
   11894: out<=0;
   11895: out<=1;
   11896: out<=0;
   11897: out<=1;
   11898: out<=1;
   11899: out<=0;
   11900: out<=0;
   11901: out<=0;
   11902: out<=0;
   11903: out<=0;
   11904: out<=1;
   11905: out<=1;
   11906: out<=0;
   11907: out<=0;
   11908: out<=1;
   11909: out<=0;
   11910: out<=1;
   11911: out<=0;
   11912: out<=1;
   11913: out<=0;
   11914: out<=0;
   11915: out<=1;
   11916: out<=1;
   11917: out<=1;
   11918: out<=1;
   11919: out<=1;
   11920: out<=1;
   11921: out<=1;
   11922: out<=0;
   11923: out<=0;
   11924: out<=1;
   11925: out<=0;
   11926: out<=1;
   11927: out<=0;
   11928: out<=1;
   11929: out<=0;
   11930: out<=0;
   11931: out<=1;
   11932: out<=1;
   11933: out<=1;
   11934: out<=1;
   11935: out<=1;
   11936: out<=1;
   11937: out<=1;
   11938: out<=0;
   11939: out<=0;
   11940: out<=1;
   11941: out<=0;
   11942: out<=1;
   11943: out<=0;
   11944: out<=1;
   11945: out<=0;
   11946: out<=0;
   11947: out<=1;
   11948: out<=1;
   11949: out<=1;
   11950: out<=1;
   11951: out<=1;
   11952: out<=1;
   11953: out<=1;
   11954: out<=0;
   11955: out<=0;
   11956: out<=1;
   11957: out<=0;
   11958: out<=1;
   11959: out<=0;
   11960: out<=1;
   11961: out<=0;
   11962: out<=0;
   11963: out<=1;
   11964: out<=1;
   11965: out<=1;
   11966: out<=1;
   11967: out<=1;
   11968: out<=1;
   11969: out<=1;
   11970: out<=0;
   11971: out<=0;
   11972: out<=1;
   11973: out<=0;
   11974: out<=1;
   11975: out<=0;
   11976: out<=1;
   11977: out<=0;
   11978: out<=0;
   11979: out<=1;
   11980: out<=1;
   11981: out<=1;
   11982: out<=1;
   11983: out<=1;
   11984: out<=0;
   11985: out<=0;
   11986: out<=1;
   11987: out<=1;
   11988: out<=0;
   11989: out<=1;
   11990: out<=0;
   11991: out<=1;
   11992: out<=0;
   11993: out<=1;
   11994: out<=1;
   11995: out<=0;
   11996: out<=0;
   11997: out<=0;
   11998: out<=0;
   11999: out<=0;
   12000: out<=0;
   12001: out<=0;
   12002: out<=1;
   12003: out<=1;
   12004: out<=0;
   12005: out<=1;
   12006: out<=0;
   12007: out<=1;
   12008: out<=0;
   12009: out<=1;
   12010: out<=1;
   12011: out<=0;
   12012: out<=0;
   12013: out<=0;
   12014: out<=0;
   12015: out<=0;
   12016: out<=1;
   12017: out<=1;
   12018: out<=0;
   12019: out<=0;
   12020: out<=1;
   12021: out<=0;
   12022: out<=1;
   12023: out<=0;
   12024: out<=1;
   12025: out<=0;
   12026: out<=0;
   12027: out<=1;
   12028: out<=1;
   12029: out<=1;
   12030: out<=1;
   12031: out<=1;
   12032: out<=1;
   12033: out<=0;
   12034: out<=1;
   12035: out<=0;
   12036: out<=0;
   12037: out<=0;
   12038: out<=1;
   12039: out<=1;
   12040: out<=0;
   12041: out<=0;
   12042: out<=0;
   12043: out<=0;
   12044: out<=1;
   12045: out<=0;
   12046: out<=0;
   12047: out<=1;
   12048: out<=1;
   12049: out<=0;
   12050: out<=1;
   12051: out<=0;
   12052: out<=0;
   12053: out<=0;
   12054: out<=1;
   12055: out<=1;
   12056: out<=0;
   12057: out<=0;
   12058: out<=0;
   12059: out<=0;
   12060: out<=1;
   12061: out<=0;
   12062: out<=0;
   12063: out<=1;
   12064: out<=0;
   12065: out<=1;
   12066: out<=0;
   12067: out<=1;
   12068: out<=1;
   12069: out<=1;
   12070: out<=0;
   12071: out<=0;
   12072: out<=1;
   12073: out<=1;
   12074: out<=1;
   12075: out<=1;
   12076: out<=0;
   12077: out<=1;
   12078: out<=1;
   12079: out<=0;
   12080: out<=0;
   12081: out<=1;
   12082: out<=0;
   12083: out<=1;
   12084: out<=1;
   12085: out<=1;
   12086: out<=0;
   12087: out<=0;
   12088: out<=1;
   12089: out<=1;
   12090: out<=1;
   12091: out<=1;
   12092: out<=0;
   12093: out<=1;
   12094: out<=1;
   12095: out<=0;
   12096: out<=1;
   12097: out<=0;
   12098: out<=1;
   12099: out<=0;
   12100: out<=0;
   12101: out<=0;
   12102: out<=1;
   12103: out<=1;
   12104: out<=0;
   12105: out<=0;
   12106: out<=0;
   12107: out<=0;
   12108: out<=1;
   12109: out<=0;
   12110: out<=0;
   12111: out<=1;
   12112: out<=0;
   12113: out<=1;
   12114: out<=0;
   12115: out<=1;
   12116: out<=1;
   12117: out<=1;
   12118: out<=0;
   12119: out<=0;
   12120: out<=1;
   12121: out<=1;
   12122: out<=1;
   12123: out<=1;
   12124: out<=0;
   12125: out<=1;
   12126: out<=1;
   12127: out<=0;
   12128: out<=1;
   12129: out<=0;
   12130: out<=1;
   12131: out<=0;
   12132: out<=0;
   12133: out<=0;
   12134: out<=1;
   12135: out<=1;
   12136: out<=0;
   12137: out<=0;
   12138: out<=0;
   12139: out<=0;
   12140: out<=1;
   12141: out<=0;
   12142: out<=0;
   12143: out<=1;
   12144: out<=0;
   12145: out<=1;
   12146: out<=0;
   12147: out<=1;
   12148: out<=1;
   12149: out<=1;
   12150: out<=0;
   12151: out<=0;
   12152: out<=1;
   12153: out<=1;
   12154: out<=1;
   12155: out<=1;
   12156: out<=0;
   12157: out<=1;
   12158: out<=1;
   12159: out<=0;
   12160: out<=1;
   12161: out<=0;
   12162: out<=1;
   12163: out<=0;
   12164: out<=0;
   12165: out<=0;
   12166: out<=1;
   12167: out<=1;
   12168: out<=0;
   12169: out<=0;
   12170: out<=0;
   12171: out<=0;
   12172: out<=1;
   12173: out<=0;
   12174: out<=0;
   12175: out<=1;
   12176: out<=0;
   12177: out<=1;
   12178: out<=0;
   12179: out<=1;
   12180: out<=1;
   12181: out<=1;
   12182: out<=0;
   12183: out<=0;
   12184: out<=1;
   12185: out<=1;
   12186: out<=1;
   12187: out<=1;
   12188: out<=0;
   12189: out<=1;
   12190: out<=1;
   12191: out<=0;
   12192: out<=0;
   12193: out<=1;
   12194: out<=0;
   12195: out<=1;
   12196: out<=1;
   12197: out<=1;
   12198: out<=0;
   12199: out<=0;
   12200: out<=1;
   12201: out<=1;
   12202: out<=1;
   12203: out<=1;
   12204: out<=0;
   12205: out<=1;
   12206: out<=1;
   12207: out<=0;
   12208: out<=1;
   12209: out<=0;
   12210: out<=1;
   12211: out<=0;
   12212: out<=0;
   12213: out<=0;
   12214: out<=1;
   12215: out<=1;
   12216: out<=0;
   12217: out<=0;
   12218: out<=0;
   12219: out<=0;
   12220: out<=1;
   12221: out<=0;
   12222: out<=0;
   12223: out<=1;
   12224: out<=1;
   12225: out<=0;
   12226: out<=1;
   12227: out<=0;
   12228: out<=0;
   12229: out<=0;
   12230: out<=1;
   12231: out<=1;
   12232: out<=0;
   12233: out<=0;
   12234: out<=0;
   12235: out<=0;
   12236: out<=1;
   12237: out<=0;
   12238: out<=0;
   12239: out<=1;
   12240: out<=1;
   12241: out<=0;
   12242: out<=1;
   12243: out<=0;
   12244: out<=0;
   12245: out<=0;
   12246: out<=1;
   12247: out<=1;
   12248: out<=0;
   12249: out<=0;
   12250: out<=0;
   12251: out<=0;
   12252: out<=1;
   12253: out<=0;
   12254: out<=0;
   12255: out<=1;
   12256: out<=1;
   12257: out<=0;
   12258: out<=1;
   12259: out<=0;
   12260: out<=0;
   12261: out<=0;
   12262: out<=1;
   12263: out<=1;
   12264: out<=0;
   12265: out<=0;
   12266: out<=0;
   12267: out<=0;
   12268: out<=1;
   12269: out<=0;
   12270: out<=0;
   12271: out<=1;
   12272: out<=1;
   12273: out<=0;
   12274: out<=1;
   12275: out<=0;
   12276: out<=0;
   12277: out<=0;
   12278: out<=1;
   12279: out<=1;
   12280: out<=0;
   12281: out<=0;
   12282: out<=0;
   12283: out<=0;
   12284: out<=1;
   12285: out<=0;
   12286: out<=0;
   12287: out<=1;
   12288: out<=0;
   12289: out<=0;
   12290: out<=1;
   12291: out<=1;
   12292: out<=1;
   12293: out<=0;
   12294: out<=1;
   12295: out<=0;
   12296: out<=0;
   12297: out<=1;
   12298: out<=1;
   12299: out<=0;
   12300: out<=1;
   12301: out<=1;
   12302: out<=1;
   12303: out<=1;
   12304: out<=1;
   12305: out<=1;
   12306: out<=0;
   12307: out<=0;
   12308: out<=0;
   12309: out<=1;
   12310: out<=0;
   12311: out<=1;
   12312: out<=1;
   12313: out<=0;
   12314: out<=0;
   12315: out<=1;
   12316: out<=0;
   12317: out<=0;
   12318: out<=0;
   12319: out<=0;
   12320: out<=1;
   12321: out<=1;
   12322: out<=0;
   12323: out<=0;
   12324: out<=0;
   12325: out<=1;
   12326: out<=0;
   12327: out<=1;
   12328: out<=1;
   12329: out<=0;
   12330: out<=0;
   12331: out<=1;
   12332: out<=0;
   12333: out<=0;
   12334: out<=0;
   12335: out<=0;
   12336: out<=0;
   12337: out<=0;
   12338: out<=1;
   12339: out<=1;
   12340: out<=1;
   12341: out<=0;
   12342: out<=1;
   12343: out<=0;
   12344: out<=0;
   12345: out<=1;
   12346: out<=1;
   12347: out<=0;
   12348: out<=1;
   12349: out<=1;
   12350: out<=1;
   12351: out<=1;
   12352: out<=1;
   12353: out<=1;
   12354: out<=0;
   12355: out<=0;
   12356: out<=0;
   12357: out<=1;
   12358: out<=0;
   12359: out<=1;
   12360: out<=1;
   12361: out<=0;
   12362: out<=0;
   12363: out<=1;
   12364: out<=0;
   12365: out<=0;
   12366: out<=0;
   12367: out<=0;
   12368: out<=1;
   12369: out<=1;
   12370: out<=0;
   12371: out<=0;
   12372: out<=0;
   12373: out<=1;
   12374: out<=0;
   12375: out<=1;
   12376: out<=1;
   12377: out<=0;
   12378: out<=0;
   12379: out<=1;
   12380: out<=0;
   12381: out<=0;
   12382: out<=0;
   12383: out<=0;
   12384: out<=1;
   12385: out<=1;
   12386: out<=0;
   12387: out<=0;
   12388: out<=0;
   12389: out<=1;
   12390: out<=0;
   12391: out<=1;
   12392: out<=1;
   12393: out<=0;
   12394: out<=0;
   12395: out<=1;
   12396: out<=0;
   12397: out<=0;
   12398: out<=0;
   12399: out<=0;
   12400: out<=1;
   12401: out<=1;
   12402: out<=0;
   12403: out<=0;
   12404: out<=0;
   12405: out<=1;
   12406: out<=0;
   12407: out<=1;
   12408: out<=1;
   12409: out<=0;
   12410: out<=0;
   12411: out<=1;
   12412: out<=0;
   12413: out<=0;
   12414: out<=0;
   12415: out<=0;
   12416: out<=1;
   12417: out<=1;
   12418: out<=0;
   12419: out<=0;
   12420: out<=0;
   12421: out<=1;
   12422: out<=0;
   12423: out<=1;
   12424: out<=1;
   12425: out<=0;
   12426: out<=0;
   12427: out<=1;
   12428: out<=0;
   12429: out<=0;
   12430: out<=0;
   12431: out<=0;
   12432: out<=1;
   12433: out<=1;
   12434: out<=0;
   12435: out<=0;
   12436: out<=0;
   12437: out<=1;
   12438: out<=0;
   12439: out<=1;
   12440: out<=1;
   12441: out<=0;
   12442: out<=0;
   12443: out<=1;
   12444: out<=0;
   12445: out<=0;
   12446: out<=0;
   12447: out<=0;
   12448: out<=0;
   12449: out<=0;
   12450: out<=1;
   12451: out<=1;
   12452: out<=1;
   12453: out<=0;
   12454: out<=1;
   12455: out<=0;
   12456: out<=0;
   12457: out<=1;
   12458: out<=1;
   12459: out<=0;
   12460: out<=1;
   12461: out<=1;
   12462: out<=1;
   12463: out<=1;
   12464: out<=0;
   12465: out<=0;
   12466: out<=1;
   12467: out<=1;
   12468: out<=1;
   12469: out<=0;
   12470: out<=1;
   12471: out<=0;
   12472: out<=0;
   12473: out<=1;
   12474: out<=1;
   12475: out<=0;
   12476: out<=1;
   12477: out<=1;
   12478: out<=1;
   12479: out<=1;
   12480: out<=0;
   12481: out<=0;
   12482: out<=1;
   12483: out<=1;
   12484: out<=1;
   12485: out<=0;
   12486: out<=1;
   12487: out<=0;
   12488: out<=0;
   12489: out<=1;
   12490: out<=1;
   12491: out<=0;
   12492: out<=1;
   12493: out<=1;
   12494: out<=1;
   12495: out<=1;
   12496: out<=1;
   12497: out<=1;
   12498: out<=0;
   12499: out<=0;
   12500: out<=0;
   12501: out<=1;
   12502: out<=0;
   12503: out<=1;
   12504: out<=1;
   12505: out<=0;
   12506: out<=0;
   12507: out<=1;
   12508: out<=0;
   12509: out<=0;
   12510: out<=0;
   12511: out<=0;
   12512: out<=0;
   12513: out<=0;
   12514: out<=1;
   12515: out<=1;
   12516: out<=1;
   12517: out<=0;
   12518: out<=1;
   12519: out<=0;
   12520: out<=0;
   12521: out<=1;
   12522: out<=1;
   12523: out<=0;
   12524: out<=1;
   12525: out<=1;
   12526: out<=1;
   12527: out<=1;
   12528: out<=1;
   12529: out<=1;
   12530: out<=0;
   12531: out<=0;
   12532: out<=0;
   12533: out<=1;
   12534: out<=0;
   12535: out<=1;
   12536: out<=1;
   12537: out<=0;
   12538: out<=0;
   12539: out<=1;
   12540: out<=0;
   12541: out<=0;
   12542: out<=0;
   12543: out<=0;
   12544: out<=0;
   12545: out<=1;
   12546: out<=0;
   12547: out<=1;
   12548: out<=0;
   12549: out<=0;
   12550: out<=1;
   12551: out<=1;
   12552: out<=1;
   12553: out<=1;
   12554: out<=1;
   12555: out<=1;
   12556: out<=1;
   12557: out<=0;
   12558: out<=0;
   12559: out<=1;
   12560: out<=0;
   12561: out<=1;
   12562: out<=0;
   12563: out<=1;
   12564: out<=0;
   12565: out<=0;
   12566: out<=1;
   12567: out<=1;
   12568: out<=1;
   12569: out<=1;
   12570: out<=1;
   12571: out<=1;
   12572: out<=1;
   12573: out<=0;
   12574: out<=0;
   12575: out<=1;
   12576: out<=0;
   12577: out<=1;
   12578: out<=0;
   12579: out<=1;
   12580: out<=0;
   12581: out<=0;
   12582: out<=1;
   12583: out<=1;
   12584: out<=1;
   12585: out<=1;
   12586: out<=1;
   12587: out<=1;
   12588: out<=1;
   12589: out<=0;
   12590: out<=0;
   12591: out<=1;
   12592: out<=0;
   12593: out<=1;
   12594: out<=0;
   12595: out<=1;
   12596: out<=0;
   12597: out<=0;
   12598: out<=1;
   12599: out<=1;
   12600: out<=1;
   12601: out<=1;
   12602: out<=1;
   12603: out<=1;
   12604: out<=1;
   12605: out<=0;
   12606: out<=0;
   12607: out<=1;
   12608: out<=1;
   12609: out<=0;
   12610: out<=1;
   12611: out<=0;
   12612: out<=1;
   12613: out<=1;
   12614: out<=0;
   12615: out<=0;
   12616: out<=0;
   12617: out<=0;
   12618: out<=0;
   12619: out<=0;
   12620: out<=0;
   12621: out<=1;
   12622: out<=1;
   12623: out<=0;
   12624: out<=0;
   12625: out<=1;
   12626: out<=0;
   12627: out<=1;
   12628: out<=0;
   12629: out<=0;
   12630: out<=1;
   12631: out<=1;
   12632: out<=1;
   12633: out<=1;
   12634: out<=1;
   12635: out<=1;
   12636: out<=1;
   12637: out<=0;
   12638: out<=0;
   12639: out<=1;
   12640: out<=0;
   12641: out<=1;
   12642: out<=0;
   12643: out<=1;
   12644: out<=0;
   12645: out<=0;
   12646: out<=1;
   12647: out<=1;
   12648: out<=1;
   12649: out<=1;
   12650: out<=1;
   12651: out<=1;
   12652: out<=1;
   12653: out<=0;
   12654: out<=0;
   12655: out<=1;
   12656: out<=1;
   12657: out<=0;
   12658: out<=1;
   12659: out<=0;
   12660: out<=1;
   12661: out<=1;
   12662: out<=0;
   12663: out<=0;
   12664: out<=0;
   12665: out<=0;
   12666: out<=0;
   12667: out<=0;
   12668: out<=0;
   12669: out<=1;
   12670: out<=1;
   12671: out<=0;
   12672: out<=1;
   12673: out<=0;
   12674: out<=1;
   12675: out<=0;
   12676: out<=1;
   12677: out<=1;
   12678: out<=0;
   12679: out<=0;
   12680: out<=0;
   12681: out<=0;
   12682: out<=0;
   12683: out<=0;
   12684: out<=0;
   12685: out<=1;
   12686: out<=1;
   12687: out<=0;
   12688: out<=0;
   12689: out<=1;
   12690: out<=0;
   12691: out<=1;
   12692: out<=0;
   12693: out<=0;
   12694: out<=1;
   12695: out<=1;
   12696: out<=1;
   12697: out<=1;
   12698: out<=1;
   12699: out<=1;
   12700: out<=1;
   12701: out<=0;
   12702: out<=0;
   12703: out<=1;
   12704: out<=1;
   12705: out<=0;
   12706: out<=1;
   12707: out<=0;
   12708: out<=1;
   12709: out<=1;
   12710: out<=0;
   12711: out<=0;
   12712: out<=0;
   12713: out<=0;
   12714: out<=0;
   12715: out<=0;
   12716: out<=0;
   12717: out<=1;
   12718: out<=1;
   12719: out<=0;
   12720: out<=0;
   12721: out<=1;
   12722: out<=0;
   12723: out<=1;
   12724: out<=0;
   12725: out<=0;
   12726: out<=1;
   12727: out<=1;
   12728: out<=1;
   12729: out<=1;
   12730: out<=1;
   12731: out<=1;
   12732: out<=1;
   12733: out<=0;
   12734: out<=0;
   12735: out<=1;
   12736: out<=0;
   12737: out<=1;
   12738: out<=0;
   12739: out<=1;
   12740: out<=0;
   12741: out<=0;
   12742: out<=1;
   12743: out<=1;
   12744: out<=1;
   12745: out<=1;
   12746: out<=1;
   12747: out<=1;
   12748: out<=1;
   12749: out<=0;
   12750: out<=0;
   12751: out<=1;
   12752: out<=0;
   12753: out<=1;
   12754: out<=0;
   12755: out<=1;
   12756: out<=0;
   12757: out<=0;
   12758: out<=1;
   12759: out<=1;
   12760: out<=1;
   12761: out<=1;
   12762: out<=1;
   12763: out<=1;
   12764: out<=1;
   12765: out<=0;
   12766: out<=0;
   12767: out<=1;
   12768: out<=1;
   12769: out<=0;
   12770: out<=1;
   12771: out<=0;
   12772: out<=1;
   12773: out<=1;
   12774: out<=0;
   12775: out<=0;
   12776: out<=0;
   12777: out<=0;
   12778: out<=0;
   12779: out<=0;
   12780: out<=0;
   12781: out<=1;
   12782: out<=1;
   12783: out<=0;
   12784: out<=1;
   12785: out<=0;
   12786: out<=1;
   12787: out<=0;
   12788: out<=1;
   12789: out<=1;
   12790: out<=0;
   12791: out<=0;
   12792: out<=0;
   12793: out<=0;
   12794: out<=0;
   12795: out<=0;
   12796: out<=0;
   12797: out<=1;
   12798: out<=1;
   12799: out<=0;
   12800: out<=0;
   12801: out<=1;
   12802: out<=1;
   12803: out<=0;
   12804: out<=0;
   12805: out<=0;
   12806: out<=0;
   12807: out<=0;
   12808: out<=0;
   12809: out<=0;
   12810: out<=1;
   12811: out<=1;
   12812: out<=0;
   12813: out<=1;
   12814: out<=0;
   12815: out<=1;
   12816: out<=0;
   12817: out<=1;
   12818: out<=1;
   12819: out<=0;
   12820: out<=0;
   12821: out<=0;
   12822: out<=0;
   12823: out<=0;
   12824: out<=0;
   12825: out<=0;
   12826: out<=1;
   12827: out<=1;
   12828: out<=0;
   12829: out<=1;
   12830: out<=0;
   12831: out<=1;
   12832: out<=1;
   12833: out<=0;
   12834: out<=0;
   12835: out<=1;
   12836: out<=1;
   12837: out<=1;
   12838: out<=1;
   12839: out<=1;
   12840: out<=1;
   12841: out<=1;
   12842: out<=0;
   12843: out<=0;
   12844: out<=1;
   12845: out<=0;
   12846: out<=1;
   12847: out<=0;
   12848: out<=1;
   12849: out<=0;
   12850: out<=0;
   12851: out<=1;
   12852: out<=1;
   12853: out<=1;
   12854: out<=1;
   12855: out<=1;
   12856: out<=1;
   12857: out<=1;
   12858: out<=0;
   12859: out<=0;
   12860: out<=1;
   12861: out<=0;
   12862: out<=1;
   12863: out<=0;
   12864: out<=1;
   12865: out<=0;
   12866: out<=0;
   12867: out<=1;
   12868: out<=1;
   12869: out<=1;
   12870: out<=1;
   12871: out<=1;
   12872: out<=1;
   12873: out<=1;
   12874: out<=0;
   12875: out<=0;
   12876: out<=1;
   12877: out<=0;
   12878: out<=1;
   12879: out<=0;
   12880: out<=0;
   12881: out<=1;
   12882: out<=1;
   12883: out<=0;
   12884: out<=0;
   12885: out<=0;
   12886: out<=0;
   12887: out<=0;
   12888: out<=0;
   12889: out<=0;
   12890: out<=1;
   12891: out<=1;
   12892: out<=0;
   12893: out<=1;
   12894: out<=0;
   12895: out<=1;
   12896: out<=1;
   12897: out<=0;
   12898: out<=0;
   12899: out<=1;
   12900: out<=1;
   12901: out<=1;
   12902: out<=1;
   12903: out<=1;
   12904: out<=1;
   12905: out<=1;
   12906: out<=0;
   12907: out<=0;
   12908: out<=1;
   12909: out<=0;
   12910: out<=1;
   12911: out<=0;
   12912: out<=0;
   12913: out<=1;
   12914: out<=1;
   12915: out<=0;
   12916: out<=0;
   12917: out<=0;
   12918: out<=0;
   12919: out<=0;
   12920: out<=0;
   12921: out<=0;
   12922: out<=1;
   12923: out<=1;
   12924: out<=0;
   12925: out<=1;
   12926: out<=0;
   12927: out<=1;
   12928: out<=1;
   12929: out<=0;
   12930: out<=0;
   12931: out<=1;
   12932: out<=1;
   12933: out<=1;
   12934: out<=1;
   12935: out<=1;
   12936: out<=1;
   12937: out<=1;
   12938: out<=0;
   12939: out<=0;
   12940: out<=1;
   12941: out<=0;
   12942: out<=1;
   12943: out<=0;
   12944: out<=0;
   12945: out<=1;
   12946: out<=1;
   12947: out<=0;
   12948: out<=0;
   12949: out<=0;
   12950: out<=0;
   12951: out<=0;
   12952: out<=0;
   12953: out<=0;
   12954: out<=1;
   12955: out<=1;
   12956: out<=0;
   12957: out<=1;
   12958: out<=0;
   12959: out<=1;
   12960: out<=0;
   12961: out<=1;
   12962: out<=1;
   12963: out<=0;
   12964: out<=0;
   12965: out<=0;
   12966: out<=0;
   12967: out<=0;
   12968: out<=0;
   12969: out<=0;
   12970: out<=1;
   12971: out<=1;
   12972: out<=0;
   12973: out<=1;
   12974: out<=0;
   12975: out<=1;
   12976: out<=1;
   12977: out<=0;
   12978: out<=0;
   12979: out<=1;
   12980: out<=1;
   12981: out<=1;
   12982: out<=1;
   12983: out<=1;
   12984: out<=1;
   12985: out<=1;
   12986: out<=0;
   12987: out<=0;
   12988: out<=1;
   12989: out<=0;
   12990: out<=1;
   12991: out<=0;
   12992: out<=0;
   12993: out<=1;
   12994: out<=1;
   12995: out<=0;
   12996: out<=0;
   12997: out<=0;
   12998: out<=0;
   12999: out<=0;
   13000: out<=0;
   13001: out<=0;
   13002: out<=1;
   13003: out<=1;
   13004: out<=0;
   13005: out<=1;
   13006: out<=0;
   13007: out<=1;
   13008: out<=0;
   13009: out<=1;
   13010: out<=1;
   13011: out<=0;
   13012: out<=0;
   13013: out<=0;
   13014: out<=0;
   13015: out<=0;
   13016: out<=0;
   13017: out<=0;
   13018: out<=1;
   13019: out<=1;
   13020: out<=0;
   13021: out<=1;
   13022: out<=0;
   13023: out<=1;
   13024: out<=0;
   13025: out<=1;
   13026: out<=1;
   13027: out<=0;
   13028: out<=0;
   13029: out<=0;
   13030: out<=0;
   13031: out<=0;
   13032: out<=0;
   13033: out<=0;
   13034: out<=1;
   13035: out<=1;
   13036: out<=0;
   13037: out<=1;
   13038: out<=0;
   13039: out<=1;
   13040: out<=0;
   13041: out<=1;
   13042: out<=1;
   13043: out<=0;
   13044: out<=0;
   13045: out<=0;
   13046: out<=0;
   13047: out<=0;
   13048: out<=0;
   13049: out<=0;
   13050: out<=1;
   13051: out<=1;
   13052: out<=0;
   13053: out<=1;
   13054: out<=0;
   13055: out<=1;
   13056: out<=0;
   13057: out<=0;
   13058: out<=0;
   13059: out<=0;
   13060: out<=1;
   13061: out<=0;
   13062: out<=0;
   13063: out<=1;
   13064: out<=1;
   13065: out<=0;
   13066: out<=1;
   13067: out<=0;
   13068: out<=0;
   13069: out<=0;
   13070: out<=1;
   13071: out<=1;
   13072: out<=1;
   13073: out<=1;
   13074: out<=1;
   13075: out<=1;
   13076: out<=0;
   13077: out<=1;
   13078: out<=1;
   13079: out<=0;
   13080: out<=0;
   13081: out<=1;
   13082: out<=0;
   13083: out<=1;
   13084: out<=1;
   13085: out<=1;
   13086: out<=0;
   13087: out<=0;
   13088: out<=0;
   13089: out<=0;
   13090: out<=0;
   13091: out<=0;
   13092: out<=1;
   13093: out<=0;
   13094: out<=0;
   13095: out<=1;
   13096: out<=1;
   13097: out<=0;
   13098: out<=1;
   13099: out<=0;
   13100: out<=0;
   13101: out<=0;
   13102: out<=1;
   13103: out<=1;
   13104: out<=1;
   13105: out<=1;
   13106: out<=1;
   13107: out<=1;
   13108: out<=0;
   13109: out<=1;
   13110: out<=1;
   13111: out<=0;
   13112: out<=0;
   13113: out<=1;
   13114: out<=0;
   13115: out<=1;
   13116: out<=1;
   13117: out<=1;
   13118: out<=0;
   13119: out<=0;
   13120: out<=1;
   13121: out<=1;
   13122: out<=1;
   13123: out<=1;
   13124: out<=0;
   13125: out<=1;
   13126: out<=1;
   13127: out<=0;
   13128: out<=0;
   13129: out<=1;
   13130: out<=0;
   13131: out<=1;
   13132: out<=1;
   13133: out<=1;
   13134: out<=0;
   13135: out<=0;
   13136: out<=1;
   13137: out<=1;
   13138: out<=1;
   13139: out<=1;
   13140: out<=0;
   13141: out<=1;
   13142: out<=1;
   13143: out<=0;
   13144: out<=0;
   13145: out<=1;
   13146: out<=0;
   13147: out<=1;
   13148: out<=1;
   13149: out<=1;
   13150: out<=0;
   13151: out<=0;
   13152: out<=0;
   13153: out<=0;
   13154: out<=0;
   13155: out<=0;
   13156: out<=1;
   13157: out<=0;
   13158: out<=0;
   13159: out<=1;
   13160: out<=1;
   13161: out<=0;
   13162: out<=1;
   13163: out<=0;
   13164: out<=0;
   13165: out<=0;
   13166: out<=1;
   13167: out<=1;
   13168: out<=0;
   13169: out<=0;
   13170: out<=0;
   13171: out<=0;
   13172: out<=1;
   13173: out<=0;
   13174: out<=0;
   13175: out<=1;
   13176: out<=1;
   13177: out<=0;
   13178: out<=1;
   13179: out<=0;
   13180: out<=0;
   13181: out<=0;
   13182: out<=1;
   13183: out<=1;
   13184: out<=1;
   13185: out<=1;
   13186: out<=1;
   13187: out<=1;
   13188: out<=0;
   13189: out<=1;
   13190: out<=1;
   13191: out<=0;
   13192: out<=0;
   13193: out<=1;
   13194: out<=0;
   13195: out<=1;
   13196: out<=1;
   13197: out<=1;
   13198: out<=0;
   13199: out<=0;
   13200: out<=1;
   13201: out<=1;
   13202: out<=1;
   13203: out<=1;
   13204: out<=0;
   13205: out<=1;
   13206: out<=1;
   13207: out<=0;
   13208: out<=0;
   13209: out<=1;
   13210: out<=0;
   13211: out<=1;
   13212: out<=1;
   13213: out<=1;
   13214: out<=0;
   13215: out<=0;
   13216: out<=1;
   13217: out<=1;
   13218: out<=1;
   13219: out<=1;
   13220: out<=0;
   13221: out<=1;
   13222: out<=1;
   13223: out<=0;
   13224: out<=0;
   13225: out<=1;
   13226: out<=0;
   13227: out<=1;
   13228: out<=1;
   13229: out<=1;
   13230: out<=0;
   13231: out<=0;
   13232: out<=1;
   13233: out<=1;
   13234: out<=1;
   13235: out<=1;
   13236: out<=0;
   13237: out<=1;
   13238: out<=1;
   13239: out<=0;
   13240: out<=0;
   13241: out<=1;
   13242: out<=0;
   13243: out<=1;
   13244: out<=1;
   13245: out<=1;
   13246: out<=0;
   13247: out<=0;
   13248: out<=0;
   13249: out<=0;
   13250: out<=0;
   13251: out<=0;
   13252: out<=1;
   13253: out<=0;
   13254: out<=0;
   13255: out<=1;
   13256: out<=1;
   13257: out<=0;
   13258: out<=1;
   13259: out<=0;
   13260: out<=0;
   13261: out<=0;
   13262: out<=1;
   13263: out<=1;
   13264: out<=1;
   13265: out<=1;
   13266: out<=1;
   13267: out<=1;
   13268: out<=0;
   13269: out<=1;
   13270: out<=1;
   13271: out<=0;
   13272: out<=0;
   13273: out<=1;
   13274: out<=0;
   13275: out<=1;
   13276: out<=1;
   13277: out<=1;
   13278: out<=0;
   13279: out<=0;
   13280: out<=1;
   13281: out<=1;
   13282: out<=1;
   13283: out<=1;
   13284: out<=0;
   13285: out<=1;
   13286: out<=1;
   13287: out<=0;
   13288: out<=0;
   13289: out<=1;
   13290: out<=0;
   13291: out<=1;
   13292: out<=1;
   13293: out<=1;
   13294: out<=0;
   13295: out<=0;
   13296: out<=0;
   13297: out<=0;
   13298: out<=0;
   13299: out<=0;
   13300: out<=1;
   13301: out<=0;
   13302: out<=0;
   13303: out<=1;
   13304: out<=1;
   13305: out<=0;
   13306: out<=1;
   13307: out<=0;
   13308: out<=0;
   13309: out<=0;
   13310: out<=1;
   13311: out<=1;
   13312: out<=0;
   13313: out<=1;
   13314: out<=0;
   13315: out<=1;
   13316: out<=1;
   13317: out<=1;
   13318: out<=0;
   13319: out<=0;
   13320: out<=0;
   13321: out<=0;
   13322: out<=0;
   13323: out<=0;
   13324: out<=1;
   13325: out<=0;
   13326: out<=0;
   13327: out<=1;
   13328: out<=1;
   13329: out<=0;
   13330: out<=1;
   13331: out<=0;
   13332: out<=0;
   13333: out<=0;
   13334: out<=1;
   13335: out<=1;
   13336: out<=1;
   13337: out<=1;
   13338: out<=1;
   13339: out<=1;
   13340: out<=0;
   13341: out<=1;
   13342: out<=1;
   13343: out<=0;
   13344: out<=1;
   13345: out<=0;
   13346: out<=1;
   13347: out<=0;
   13348: out<=0;
   13349: out<=0;
   13350: out<=1;
   13351: out<=1;
   13352: out<=1;
   13353: out<=1;
   13354: out<=1;
   13355: out<=1;
   13356: out<=0;
   13357: out<=1;
   13358: out<=1;
   13359: out<=0;
   13360: out<=0;
   13361: out<=1;
   13362: out<=0;
   13363: out<=1;
   13364: out<=1;
   13365: out<=1;
   13366: out<=0;
   13367: out<=0;
   13368: out<=0;
   13369: out<=0;
   13370: out<=0;
   13371: out<=0;
   13372: out<=1;
   13373: out<=0;
   13374: out<=0;
   13375: out<=1;
   13376: out<=1;
   13377: out<=0;
   13378: out<=1;
   13379: out<=0;
   13380: out<=0;
   13381: out<=0;
   13382: out<=1;
   13383: out<=1;
   13384: out<=1;
   13385: out<=1;
   13386: out<=1;
   13387: out<=1;
   13388: out<=0;
   13389: out<=1;
   13390: out<=1;
   13391: out<=0;
   13392: out<=1;
   13393: out<=0;
   13394: out<=1;
   13395: out<=0;
   13396: out<=0;
   13397: out<=0;
   13398: out<=1;
   13399: out<=1;
   13400: out<=1;
   13401: out<=1;
   13402: out<=1;
   13403: out<=1;
   13404: out<=0;
   13405: out<=1;
   13406: out<=1;
   13407: out<=0;
   13408: out<=1;
   13409: out<=0;
   13410: out<=1;
   13411: out<=0;
   13412: out<=0;
   13413: out<=0;
   13414: out<=1;
   13415: out<=1;
   13416: out<=1;
   13417: out<=1;
   13418: out<=1;
   13419: out<=1;
   13420: out<=0;
   13421: out<=1;
   13422: out<=1;
   13423: out<=0;
   13424: out<=1;
   13425: out<=0;
   13426: out<=1;
   13427: out<=0;
   13428: out<=0;
   13429: out<=0;
   13430: out<=1;
   13431: out<=1;
   13432: out<=1;
   13433: out<=1;
   13434: out<=1;
   13435: out<=1;
   13436: out<=0;
   13437: out<=1;
   13438: out<=1;
   13439: out<=0;
   13440: out<=1;
   13441: out<=0;
   13442: out<=1;
   13443: out<=0;
   13444: out<=0;
   13445: out<=0;
   13446: out<=1;
   13447: out<=1;
   13448: out<=1;
   13449: out<=1;
   13450: out<=1;
   13451: out<=1;
   13452: out<=0;
   13453: out<=1;
   13454: out<=1;
   13455: out<=0;
   13456: out<=1;
   13457: out<=0;
   13458: out<=1;
   13459: out<=0;
   13460: out<=0;
   13461: out<=0;
   13462: out<=1;
   13463: out<=1;
   13464: out<=1;
   13465: out<=1;
   13466: out<=1;
   13467: out<=1;
   13468: out<=0;
   13469: out<=1;
   13470: out<=1;
   13471: out<=0;
   13472: out<=0;
   13473: out<=1;
   13474: out<=0;
   13475: out<=1;
   13476: out<=1;
   13477: out<=1;
   13478: out<=0;
   13479: out<=0;
   13480: out<=0;
   13481: out<=0;
   13482: out<=0;
   13483: out<=0;
   13484: out<=1;
   13485: out<=0;
   13486: out<=0;
   13487: out<=1;
   13488: out<=0;
   13489: out<=1;
   13490: out<=0;
   13491: out<=1;
   13492: out<=1;
   13493: out<=1;
   13494: out<=0;
   13495: out<=0;
   13496: out<=0;
   13497: out<=0;
   13498: out<=0;
   13499: out<=0;
   13500: out<=1;
   13501: out<=0;
   13502: out<=0;
   13503: out<=1;
   13504: out<=0;
   13505: out<=1;
   13506: out<=0;
   13507: out<=1;
   13508: out<=1;
   13509: out<=1;
   13510: out<=0;
   13511: out<=0;
   13512: out<=0;
   13513: out<=0;
   13514: out<=0;
   13515: out<=0;
   13516: out<=1;
   13517: out<=0;
   13518: out<=0;
   13519: out<=1;
   13520: out<=1;
   13521: out<=0;
   13522: out<=1;
   13523: out<=0;
   13524: out<=0;
   13525: out<=0;
   13526: out<=1;
   13527: out<=1;
   13528: out<=1;
   13529: out<=1;
   13530: out<=1;
   13531: out<=1;
   13532: out<=0;
   13533: out<=1;
   13534: out<=1;
   13535: out<=0;
   13536: out<=0;
   13537: out<=1;
   13538: out<=0;
   13539: out<=1;
   13540: out<=1;
   13541: out<=1;
   13542: out<=0;
   13543: out<=0;
   13544: out<=0;
   13545: out<=0;
   13546: out<=0;
   13547: out<=0;
   13548: out<=1;
   13549: out<=0;
   13550: out<=0;
   13551: out<=1;
   13552: out<=1;
   13553: out<=0;
   13554: out<=1;
   13555: out<=0;
   13556: out<=0;
   13557: out<=0;
   13558: out<=1;
   13559: out<=1;
   13560: out<=1;
   13561: out<=1;
   13562: out<=1;
   13563: out<=1;
   13564: out<=0;
   13565: out<=1;
   13566: out<=1;
   13567: out<=0;
   13568: out<=1;
   13569: out<=1;
   13570: out<=0;
   13571: out<=0;
   13572: out<=1;
   13573: out<=0;
   13574: out<=1;
   13575: out<=0;
   13576: out<=0;
   13577: out<=1;
   13578: out<=1;
   13579: out<=0;
   13580: out<=0;
   13581: out<=0;
   13582: out<=0;
   13583: out<=0;
   13584: out<=1;
   13585: out<=1;
   13586: out<=0;
   13587: out<=0;
   13588: out<=1;
   13589: out<=0;
   13590: out<=1;
   13591: out<=0;
   13592: out<=0;
   13593: out<=1;
   13594: out<=1;
   13595: out<=0;
   13596: out<=0;
   13597: out<=0;
   13598: out<=0;
   13599: out<=0;
   13600: out<=1;
   13601: out<=1;
   13602: out<=0;
   13603: out<=0;
   13604: out<=1;
   13605: out<=0;
   13606: out<=1;
   13607: out<=0;
   13608: out<=0;
   13609: out<=1;
   13610: out<=1;
   13611: out<=0;
   13612: out<=0;
   13613: out<=0;
   13614: out<=0;
   13615: out<=0;
   13616: out<=1;
   13617: out<=1;
   13618: out<=0;
   13619: out<=0;
   13620: out<=1;
   13621: out<=0;
   13622: out<=1;
   13623: out<=0;
   13624: out<=0;
   13625: out<=1;
   13626: out<=1;
   13627: out<=0;
   13628: out<=0;
   13629: out<=0;
   13630: out<=0;
   13631: out<=0;
   13632: out<=0;
   13633: out<=0;
   13634: out<=1;
   13635: out<=1;
   13636: out<=0;
   13637: out<=1;
   13638: out<=0;
   13639: out<=1;
   13640: out<=1;
   13641: out<=0;
   13642: out<=0;
   13643: out<=1;
   13644: out<=1;
   13645: out<=1;
   13646: out<=1;
   13647: out<=1;
   13648: out<=1;
   13649: out<=1;
   13650: out<=0;
   13651: out<=0;
   13652: out<=1;
   13653: out<=0;
   13654: out<=1;
   13655: out<=0;
   13656: out<=0;
   13657: out<=1;
   13658: out<=1;
   13659: out<=0;
   13660: out<=0;
   13661: out<=0;
   13662: out<=0;
   13663: out<=0;
   13664: out<=1;
   13665: out<=1;
   13666: out<=0;
   13667: out<=0;
   13668: out<=1;
   13669: out<=0;
   13670: out<=1;
   13671: out<=0;
   13672: out<=0;
   13673: out<=1;
   13674: out<=1;
   13675: out<=0;
   13676: out<=0;
   13677: out<=0;
   13678: out<=0;
   13679: out<=0;
   13680: out<=0;
   13681: out<=0;
   13682: out<=1;
   13683: out<=1;
   13684: out<=0;
   13685: out<=1;
   13686: out<=0;
   13687: out<=1;
   13688: out<=1;
   13689: out<=0;
   13690: out<=0;
   13691: out<=1;
   13692: out<=1;
   13693: out<=1;
   13694: out<=1;
   13695: out<=1;
   13696: out<=0;
   13697: out<=0;
   13698: out<=1;
   13699: out<=1;
   13700: out<=0;
   13701: out<=1;
   13702: out<=0;
   13703: out<=1;
   13704: out<=1;
   13705: out<=0;
   13706: out<=0;
   13707: out<=1;
   13708: out<=1;
   13709: out<=1;
   13710: out<=1;
   13711: out<=1;
   13712: out<=1;
   13713: out<=1;
   13714: out<=0;
   13715: out<=0;
   13716: out<=1;
   13717: out<=0;
   13718: out<=1;
   13719: out<=0;
   13720: out<=0;
   13721: out<=1;
   13722: out<=1;
   13723: out<=0;
   13724: out<=0;
   13725: out<=0;
   13726: out<=0;
   13727: out<=0;
   13728: out<=0;
   13729: out<=0;
   13730: out<=1;
   13731: out<=1;
   13732: out<=0;
   13733: out<=1;
   13734: out<=0;
   13735: out<=1;
   13736: out<=1;
   13737: out<=0;
   13738: out<=0;
   13739: out<=1;
   13740: out<=1;
   13741: out<=1;
   13742: out<=1;
   13743: out<=1;
   13744: out<=1;
   13745: out<=1;
   13746: out<=0;
   13747: out<=0;
   13748: out<=1;
   13749: out<=0;
   13750: out<=1;
   13751: out<=0;
   13752: out<=0;
   13753: out<=1;
   13754: out<=1;
   13755: out<=0;
   13756: out<=0;
   13757: out<=0;
   13758: out<=0;
   13759: out<=0;
   13760: out<=1;
   13761: out<=1;
   13762: out<=0;
   13763: out<=0;
   13764: out<=1;
   13765: out<=0;
   13766: out<=1;
   13767: out<=0;
   13768: out<=0;
   13769: out<=1;
   13770: out<=1;
   13771: out<=0;
   13772: out<=0;
   13773: out<=0;
   13774: out<=0;
   13775: out<=0;
   13776: out<=1;
   13777: out<=1;
   13778: out<=0;
   13779: out<=0;
   13780: out<=1;
   13781: out<=0;
   13782: out<=1;
   13783: out<=0;
   13784: out<=0;
   13785: out<=1;
   13786: out<=1;
   13787: out<=0;
   13788: out<=0;
   13789: out<=0;
   13790: out<=0;
   13791: out<=0;
   13792: out<=0;
   13793: out<=0;
   13794: out<=1;
   13795: out<=1;
   13796: out<=0;
   13797: out<=1;
   13798: out<=0;
   13799: out<=1;
   13800: out<=1;
   13801: out<=0;
   13802: out<=0;
   13803: out<=1;
   13804: out<=1;
   13805: out<=1;
   13806: out<=1;
   13807: out<=1;
   13808: out<=0;
   13809: out<=0;
   13810: out<=1;
   13811: out<=1;
   13812: out<=0;
   13813: out<=1;
   13814: out<=0;
   13815: out<=1;
   13816: out<=1;
   13817: out<=0;
   13818: out<=0;
   13819: out<=1;
   13820: out<=1;
   13821: out<=1;
   13822: out<=1;
   13823: out<=1;
   13824: out<=1;
   13825: out<=1;
   13826: out<=1;
   13827: out<=1;
   13828: out<=1;
   13829: out<=0;
   13830: out<=0;
   13831: out<=1;
   13832: out<=1;
   13833: out<=0;
   13834: out<=1;
   13835: out<=0;
   13836: out<=1;
   13837: out<=1;
   13838: out<=0;
   13839: out<=0;
   13840: out<=1;
   13841: out<=1;
   13842: out<=1;
   13843: out<=1;
   13844: out<=1;
   13845: out<=0;
   13846: out<=0;
   13847: out<=1;
   13848: out<=1;
   13849: out<=0;
   13850: out<=1;
   13851: out<=0;
   13852: out<=1;
   13853: out<=1;
   13854: out<=0;
   13855: out<=0;
   13856: out<=0;
   13857: out<=0;
   13858: out<=0;
   13859: out<=0;
   13860: out<=0;
   13861: out<=1;
   13862: out<=1;
   13863: out<=0;
   13864: out<=0;
   13865: out<=1;
   13866: out<=0;
   13867: out<=1;
   13868: out<=0;
   13869: out<=0;
   13870: out<=1;
   13871: out<=1;
   13872: out<=0;
   13873: out<=0;
   13874: out<=0;
   13875: out<=0;
   13876: out<=0;
   13877: out<=1;
   13878: out<=1;
   13879: out<=0;
   13880: out<=0;
   13881: out<=1;
   13882: out<=0;
   13883: out<=1;
   13884: out<=0;
   13885: out<=0;
   13886: out<=1;
   13887: out<=1;
   13888: out<=0;
   13889: out<=0;
   13890: out<=0;
   13891: out<=0;
   13892: out<=0;
   13893: out<=1;
   13894: out<=1;
   13895: out<=0;
   13896: out<=0;
   13897: out<=1;
   13898: out<=0;
   13899: out<=1;
   13900: out<=0;
   13901: out<=0;
   13902: out<=1;
   13903: out<=1;
   13904: out<=1;
   13905: out<=1;
   13906: out<=1;
   13907: out<=1;
   13908: out<=1;
   13909: out<=0;
   13910: out<=0;
   13911: out<=1;
   13912: out<=1;
   13913: out<=0;
   13914: out<=1;
   13915: out<=0;
   13916: out<=1;
   13917: out<=1;
   13918: out<=0;
   13919: out<=0;
   13920: out<=0;
   13921: out<=0;
   13922: out<=0;
   13923: out<=0;
   13924: out<=0;
   13925: out<=1;
   13926: out<=1;
   13927: out<=0;
   13928: out<=0;
   13929: out<=1;
   13930: out<=0;
   13931: out<=1;
   13932: out<=0;
   13933: out<=0;
   13934: out<=1;
   13935: out<=1;
   13936: out<=1;
   13937: out<=1;
   13938: out<=1;
   13939: out<=1;
   13940: out<=1;
   13941: out<=0;
   13942: out<=0;
   13943: out<=1;
   13944: out<=1;
   13945: out<=0;
   13946: out<=1;
   13947: out<=0;
   13948: out<=1;
   13949: out<=1;
   13950: out<=0;
   13951: out<=0;
   13952: out<=0;
   13953: out<=0;
   13954: out<=0;
   13955: out<=0;
   13956: out<=0;
   13957: out<=1;
   13958: out<=1;
   13959: out<=0;
   13960: out<=0;
   13961: out<=1;
   13962: out<=0;
   13963: out<=1;
   13964: out<=0;
   13965: out<=0;
   13966: out<=1;
   13967: out<=1;
   13968: out<=1;
   13969: out<=1;
   13970: out<=1;
   13971: out<=1;
   13972: out<=1;
   13973: out<=0;
   13974: out<=0;
   13975: out<=1;
   13976: out<=1;
   13977: out<=0;
   13978: out<=1;
   13979: out<=0;
   13980: out<=1;
   13981: out<=1;
   13982: out<=0;
   13983: out<=0;
   13984: out<=1;
   13985: out<=1;
   13986: out<=1;
   13987: out<=1;
   13988: out<=1;
   13989: out<=0;
   13990: out<=0;
   13991: out<=1;
   13992: out<=1;
   13993: out<=0;
   13994: out<=1;
   13995: out<=0;
   13996: out<=1;
   13997: out<=1;
   13998: out<=0;
   13999: out<=0;
   14000: out<=0;
   14001: out<=0;
   14002: out<=0;
   14003: out<=0;
   14004: out<=0;
   14005: out<=1;
   14006: out<=1;
   14007: out<=0;
   14008: out<=0;
   14009: out<=1;
   14010: out<=0;
   14011: out<=1;
   14012: out<=0;
   14013: out<=0;
   14014: out<=1;
   14015: out<=1;
   14016: out<=1;
   14017: out<=1;
   14018: out<=1;
   14019: out<=1;
   14020: out<=1;
   14021: out<=0;
   14022: out<=0;
   14023: out<=1;
   14024: out<=1;
   14025: out<=0;
   14026: out<=1;
   14027: out<=0;
   14028: out<=1;
   14029: out<=1;
   14030: out<=0;
   14031: out<=0;
   14032: out<=1;
   14033: out<=1;
   14034: out<=1;
   14035: out<=1;
   14036: out<=1;
   14037: out<=0;
   14038: out<=0;
   14039: out<=1;
   14040: out<=1;
   14041: out<=0;
   14042: out<=1;
   14043: out<=0;
   14044: out<=1;
   14045: out<=1;
   14046: out<=0;
   14047: out<=0;
   14048: out<=1;
   14049: out<=1;
   14050: out<=1;
   14051: out<=1;
   14052: out<=1;
   14053: out<=0;
   14054: out<=0;
   14055: out<=1;
   14056: out<=1;
   14057: out<=0;
   14058: out<=1;
   14059: out<=0;
   14060: out<=1;
   14061: out<=1;
   14062: out<=0;
   14063: out<=0;
   14064: out<=1;
   14065: out<=1;
   14066: out<=1;
   14067: out<=1;
   14068: out<=1;
   14069: out<=0;
   14070: out<=0;
   14071: out<=1;
   14072: out<=1;
   14073: out<=0;
   14074: out<=1;
   14075: out<=0;
   14076: out<=1;
   14077: out<=1;
   14078: out<=0;
   14079: out<=0;
   14080: out<=0;
   14081: out<=1;
   14082: out<=1;
   14083: out<=0;
   14084: out<=1;
   14085: out<=1;
   14086: out<=1;
   14087: out<=1;
   14088: out<=1;
   14089: out<=1;
   14090: out<=0;
   14091: out<=0;
   14092: out<=0;
   14093: out<=1;
   14094: out<=0;
   14095: out<=1;
   14096: out<=1;
   14097: out<=0;
   14098: out<=0;
   14099: out<=1;
   14100: out<=0;
   14101: out<=0;
   14102: out<=0;
   14103: out<=0;
   14104: out<=0;
   14105: out<=0;
   14106: out<=1;
   14107: out<=1;
   14108: out<=1;
   14109: out<=0;
   14110: out<=1;
   14111: out<=0;
   14112: out<=0;
   14113: out<=1;
   14114: out<=1;
   14115: out<=0;
   14116: out<=1;
   14117: out<=1;
   14118: out<=1;
   14119: out<=1;
   14120: out<=1;
   14121: out<=1;
   14122: out<=0;
   14123: out<=0;
   14124: out<=0;
   14125: out<=1;
   14126: out<=0;
   14127: out<=1;
   14128: out<=1;
   14129: out<=0;
   14130: out<=0;
   14131: out<=1;
   14132: out<=0;
   14133: out<=0;
   14134: out<=0;
   14135: out<=0;
   14136: out<=0;
   14137: out<=0;
   14138: out<=1;
   14139: out<=1;
   14140: out<=1;
   14141: out<=0;
   14142: out<=1;
   14143: out<=0;
   14144: out<=1;
   14145: out<=0;
   14146: out<=0;
   14147: out<=1;
   14148: out<=0;
   14149: out<=0;
   14150: out<=0;
   14151: out<=0;
   14152: out<=0;
   14153: out<=0;
   14154: out<=1;
   14155: out<=1;
   14156: out<=1;
   14157: out<=0;
   14158: out<=1;
   14159: out<=0;
   14160: out<=1;
   14161: out<=0;
   14162: out<=0;
   14163: out<=1;
   14164: out<=0;
   14165: out<=0;
   14166: out<=0;
   14167: out<=0;
   14168: out<=0;
   14169: out<=0;
   14170: out<=1;
   14171: out<=1;
   14172: out<=1;
   14173: out<=0;
   14174: out<=1;
   14175: out<=0;
   14176: out<=0;
   14177: out<=1;
   14178: out<=1;
   14179: out<=0;
   14180: out<=1;
   14181: out<=1;
   14182: out<=1;
   14183: out<=1;
   14184: out<=1;
   14185: out<=1;
   14186: out<=0;
   14187: out<=0;
   14188: out<=0;
   14189: out<=1;
   14190: out<=0;
   14191: out<=1;
   14192: out<=0;
   14193: out<=1;
   14194: out<=1;
   14195: out<=0;
   14196: out<=1;
   14197: out<=1;
   14198: out<=1;
   14199: out<=1;
   14200: out<=1;
   14201: out<=1;
   14202: out<=0;
   14203: out<=0;
   14204: out<=0;
   14205: out<=1;
   14206: out<=0;
   14207: out<=1;
   14208: out<=1;
   14209: out<=0;
   14210: out<=0;
   14211: out<=1;
   14212: out<=0;
   14213: out<=0;
   14214: out<=0;
   14215: out<=0;
   14216: out<=0;
   14217: out<=0;
   14218: out<=1;
   14219: out<=1;
   14220: out<=1;
   14221: out<=0;
   14222: out<=1;
   14223: out<=0;
   14224: out<=1;
   14225: out<=0;
   14226: out<=0;
   14227: out<=1;
   14228: out<=0;
   14229: out<=0;
   14230: out<=0;
   14231: out<=0;
   14232: out<=0;
   14233: out<=0;
   14234: out<=1;
   14235: out<=1;
   14236: out<=1;
   14237: out<=0;
   14238: out<=1;
   14239: out<=0;
   14240: out<=1;
   14241: out<=0;
   14242: out<=0;
   14243: out<=1;
   14244: out<=0;
   14245: out<=0;
   14246: out<=0;
   14247: out<=0;
   14248: out<=0;
   14249: out<=0;
   14250: out<=1;
   14251: out<=1;
   14252: out<=1;
   14253: out<=0;
   14254: out<=1;
   14255: out<=0;
   14256: out<=1;
   14257: out<=0;
   14258: out<=0;
   14259: out<=1;
   14260: out<=0;
   14261: out<=0;
   14262: out<=0;
   14263: out<=0;
   14264: out<=0;
   14265: out<=0;
   14266: out<=1;
   14267: out<=1;
   14268: out<=1;
   14269: out<=0;
   14270: out<=1;
   14271: out<=0;
   14272: out<=0;
   14273: out<=1;
   14274: out<=1;
   14275: out<=0;
   14276: out<=1;
   14277: out<=1;
   14278: out<=1;
   14279: out<=1;
   14280: out<=1;
   14281: out<=1;
   14282: out<=0;
   14283: out<=0;
   14284: out<=0;
   14285: out<=1;
   14286: out<=0;
   14287: out<=1;
   14288: out<=1;
   14289: out<=0;
   14290: out<=0;
   14291: out<=1;
   14292: out<=0;
   14293: out<=0;
   14294: out<=0;
   14295: out<=0;
   14296: out<=0;
   14297: out<=0;
   14298: out<=1;
   14299: out<=1;
   14300: out<=1;
   14301: out<=0;
   14302: out<=1;
   14303: out<=0;
   14304: out<=1;
   14305: out<=0;
   14306: out<=0;
   14307: out<=1;
   14308: out<=0;
   14309: out<=0;
   14310: out<=0;
   14311: out<=0;
   14312: out<=0;
   14313: out<=0;
   14314: out<=1;
   14315: out<=1;
   14316: out<=1;
   14317: out<=0;
   14318: out<=1;
   14319: out<=0;
   14320: out<=0;
   14321: out<=1;
   14322: out<=1;
   14323: out<=0;
   14324: out<=1;
   14325: out<=1;
   14326: out<=1;
   14327: out<=1;
   14328: out<=1;
   14329: out<=1;
   14330: out<=0;
   14331: out<=0;
   14332: out<=0;
   14333: out<=1;
   14334: out<=0;
   14335: out<=1;
   14336: out<=0;
   14337: out<=1;
   14338: out<=1;
   14339: out<=0;
   14340: out<=1;
   14341: out<=1;
   14342: out<=1;
   14343: out<=1;
   14344: out<=0;
   14345: out<=0;
   14346: out<=1;
   14347: out<=1;
   14348: out<=1;
   14349: out<=0;
   14350: out<=1;
   14351: out<=0;
   14352: out<=1;
   14353: out<=0;
   14354: out<=0;
   14355: out<=1;
   14356: out<=0;
   14357: out<=0;
   14358: out<=0;
   14359: out<=0;
   14360: out<=1;
   14361: out<=1;
   14362: out<=0;
   14363: out<=0;
   14364: out<=0;
   14365: out<=1;
   14366: out<=0;
   14367: out<=1;
   14368: out<=1;
   14369: out<=0;
   14370: out<=0;
   14371: out<=1;
   14372: out<=0;
   14373: out<=0;
   14374: out<=0;
   14375: out<=0;
   14376: out<=1;
   14377: out<=1;
   14378: out<=0;
   14379: out<=0;
   14380: out<=0;
   14381: out<=1;
   14382: out<=0;
   14383: out<=1;
   14384: out<=0;
   14385: out<=1;
   14386: out<=1;
   14387: out<=0;
   14388: out<=1;
   14389: out<=1;
   14390: out<=1;
   14391: out<=1;
   14392: out<=0;
   14393: out<=0;
   14394: out<=1;
   14395: out<=1;
   14396: out<=1;
   14397: out<=0;
   14398: out<=1;
   14399: out<=0;
   14400: out<=1;
   14401: out<=0;
   14402: out<=0;
   14403: out<=1;
   14404: out<=0;
   14405: out<=0;
   14406: out<=0;
   14407: out<=0;
   14408: out<=1;
   14409: out<=1;
   14410: out<=0;
   14411: out<=0;
   14412: out<=0;
   14413: out<=1;
   14414: out<=0;
   14415: out<=1;
   14416: out<=1;
   14417: out<=0;
   14418: out<=0;
   14419: out<=1;
   14420: out<=0;
   14421: out<=0;
   14422: out<=0;
   14423: out<=0;
   14424: out<=1;
   14425: out<=1;
   14426: out<=0;
   14427: out<=0;
   14428: out<=0;
   14429: out<=1;
   14430: out<=0;
   14431: out<=1;
   14432: out<=1;
   14433: out<=0;
   14434: out<=0;
   14435: out<=1;
   14436: out<=0;
   14437: out<=0;
   14438: out<=0;
   14439: out<=0;
   14440: out<=1;
   14441: out<=1;
   14442: out<=0;
   14443: out<=0;
   14444: out<=0;
   14445: out<=1;
   14446: out<=0;
   14447: out<=1;
   14448: out<=1;
   14449: out<=0;
   14450: out<=0;
   14451: out<=1;
   14452: out<=0;
   14453: out<=0;
   14454: out<=0;
   14455: out<=0;
   14456: out<=1;
   14457: out<=1;
   14458: out<=0;
   14459: out<=0;
   14460: out<=0;
   14461: out<=1;
   14462: out<=0;
   14463: out<=1;
   14464: out<=1;
   14465: out<=0;
   14466: out<=0;
   14467: out<=1;
   14468: out<=0;
   14469: out<=0;
   14470: out<=0;
   14471: out<=0;
   14472: out<=1;
   14473: out<=1;
   14474: out<=0;
   14475: out<=0;
   14476: out<=0;
   14477: out<=1;
   14478: out<=0;
   14479: out<=1;
   14480: out<=1;
   14481: out<=0;
   14482: out<=0;
   14483: out<=1;
   14484: out<=0;
   14485: out<=0;
   14486: out<=0;
   14487: out<=0;
   14488: out<=1;
   14489: out<=1;
   14490: out<=0;
   14491: out<=0;
   14492: out<=0;
   14493: out<=1;
   14494: out<=0;
   14495: out<=1;
   14496: out<=0;
   14497: out<=1;
   14498: out<=1;
   14499: out<=0;
   14500: out<=1;
   14501: out<=1;
   14502: out<=1;
   14503: out<=1;
   14504: out<=0;
   14505: out<=0;
   14506: out<=1;
   14507: out<=1;
   14508: out<=1;
   14509: out<=0;
   14510: out<=1;
   14511: out<=0;
   14512: out<=0;
   14513: out<=1;
   14514: out<=1;
   14515: out<=0;
   14516: out<=1;
   14517: out<=1;
   14518: out<=1;
   14519: out<=1;
   14520: out<=0;
   14521: out<=0;
   14522: out<=1;
   14523: out<=1;
   14524: out<=1;
   14525: out<=0;
   14526: out<=1;
   14527: out<=0;
   14528: out<=0;
   14529: out<=1;
   14530: out<=1;
   14531: out<=0;
   14532: out<=1;
   14533: out<=1;
   14534: out<=1;
   14535: out<=1;
   14536: out<=0;
   14537: out<=0;
   14538: out<=1;
   14539: out<=1;
   14540: out<=1;
   14541: out<=0;
   14542: out<=1;
   14543: out<=0;
   14544: out<=1;
   14545: out<=0;
   14546: out<=0;
   14547: out<=1;
   14548: out<=0;
   14549: out<=0;
   14550: out<=0;
   14551: out<=0;
   14552: out<=1;
   14553: out<=1;
   14554: out<=0;
   14555: out<=0;
   14556: out<=0;
   14557: out<=1;
   14558: out<=0;
   14559: out<=1;
   14560: out<=0;
   14561: out<=1;
   14562: out<=1;
   14563: out<=0;
   14564: out<=1;
   14565: out<=1;
   14566: out<=1;
   14567: out<=1;
   14568: out<=0;
   14569: out<=0;
   14570: out<=1;
   14571: out<=1;
   14572: out<=1;
   14573: out<=0;
   14574: out<=1;
   14575: out<=0;
   14576: out<=1;
   14577: out<=0;
   14578: out<=0;
   14579: out<=1;
   14580: out<=0;
   14581: out<=0;
   14582: out<=0;
   14583: out<=0;
   14584: out<=1;
   14585: out<=1;
   14586: out<=0;
   14587: out<=0;
   14588: out<=0;
   14589: out<=1;
   14590: out<=0;
   14591: out<=1;
   14592: out<=1;
   14593: out<=1;
   14594: out<=1;
   14595: out<=1;
   14596: out<=1;
   14597: out<=0;
   14598: out<=0;
   14599: out<=1;
   14600: out<=0;
   14601: out<=1;
   14602: out<=0;
   14603: out<=1;
   14604: out<=0;
   14605: out<=0;
   14606: out<=1;
   14607: out<=1;
   14608: out<=1;
   14609: out<=1;
   14610: out<=1;
   14611: out<=1;
   14612: out<=1;
   14613: out<=0;
   14614: out<=0;
   14615: out<=1;
   14616: out<=0;
   14617: out<=1;
   14618: out<=0;
   14619: out<=1;
   14620: out<=0;
   14621: out<=0;
   14622: out<=1;
   14623: out<=1;
   14624: out<=1;
   14625: out<=1;
   14626: out<=1;
   14627: out<=1;
   14628: out<=1;
   14629: out<=0;
   14630: out<=0;
   14631: out<=1;
   14632: out<=0;
   14633: out<=1;
   14634: out<=0;
   14635: out<=1;
   14636: out<=0;
   14637: out<=0;
   14638: out<=1;
   14639: out<=1;
   14640: out<=1;
   14641: out<=1;
   14642: out<=1;
   14643: out<=1;
   14644: out<=1;
   14645: out<=0;
   14646: out<=0;
   14647: out<=1;
   14648: out<=0;
   14649: out<=1;
   14650: out<=0;
   14651: out<=1;
   14652: out<=0;
   14653: out<=0;
   14654: out<=1;
   14655: out<=1;
   14656: out<=0;
   14657: out<=0;
   14658: out<=0;
   14659: out<=0;
   14660: out<=0;
   14661: out<=1;
   14662: out<=1;
   14663: out<=0;
   14664: out<=1;
   14665: out<=0;
   14666: out<=1;
   14667: out<=0;
   14668: out<=1;
   14669: out<=1;
   14670: out<=0;
   14671: out<=0;
   14672: out<=1;
   14673: out<=1;
   14674: out<=1;
   14675: out<=1;
   14676: out<=1;
   14677: out<=0;
   14678: out<=0;
   14679: out<=1;
   14680: out<=0;
   14681: out<=1;
   14682: out<=0;
   14683: out<=1;
   14684: out<=0;
   14685: out<=0;
   14686: out<=1;
   14687: out<=1;
   14688: out<=1;
   14689: out<=1;
   14690: out<=1;
   14691: out<=1;
   14692: out<=1;
   14693: out<=0;
   14694: out<=0;
   14695: out<=1;
   14696: out<=0;
   14697: out<=1;
   14698: out<=0;
   14699: out<=1;
   14700: out<=0;
   14701: out<=0;
   14702: out<=1;
   14703: out<=1;
   14704: out<=0;
   14705: out<=0;
   14706: out<=0;
   14707: out<=0;
   14708: out<=0;
   14709: out<=1;
   14710: out<=1;
   14711: out<=0;
   14712: out<=1;
   14713: out<=0;
   14714: out<=1;
   14715: out<=0;
   14716: out<=1;
   14717: out<=1;
   14718: out<=0;
   14719: out<=0;
   14720: out<=0;
   14721: out<=0;
   14722: out<=0;
   14723: out<=0;
   14724: out<=0;
   14725: out<=1;
   14726: out<=1;
   14727: out<=0;
   14728: out<=1;
   14729: out<=0;
   14730: out<=1;
   14731: out<=0;
   14732: out<=1;
   14733: out<=1;
   14734: out<=0;
   14735: out<=0;
   14736: out<=1;
   14737: out<=1;
   14738: out<=1;
   14739: out<=1;
   14740: out<=1;
   14741: out<=0;
   14742: out<=0;
   14743: out<=1;
   14744: out<=0;
   14745: out<=1;
   14746: out<=0;
   14747: out<=1;
   14748: out<=0;
   14749: out<=0;
   14750: out<=1;
   14751: out<=1;
   14752: out<=0;
   14753: out<=0;
   14754: out<=0;
   14755: out<=0;
   14756: out<=0;
   14757: out<=1;
   14758: out<=1;
   14759: out<=0;
   14760: out<=1;
   14761: out<=0;
   14762: out<=1;
   14763: out<=0;
   14764: out<=1;
   14765: out<=1;
   14766: out<=0;
   14767: out<=0;
   14768: out<=1;
   14769: out<=1;
   14770: out<=1;
   14771: out<=1;
   14772: out<=1;
   14773: out<=0;
   14774: out<=0;
   14775: out<=1;
   14776: out<=0;
   14777: out<=1;
   14778: out<=0;
   14779: out<=1;
   14780: out<=0;
   14781: out<=0;
   14782: out<=1;
   14783: out<=1;
   14784: out<=1;
   14785: out<=1;
   14786: out<=1;
   14787: out<=1;
   14788: out<=1;
   14789: out<=0;
   14790: out<=0;
   14791: out<=1;
   14792: out<=0;
   14793: out<=1;
   14794: out<=0;
   14795: out<=1;
   14796: out<=0;
   14797: out<=0;
   14798: out<=1;
   14799: out<=1;
   14800: out<=1;
   14801: out<=1;
   14802: out<=1;
   14803: out<=1;
   14804: out<=1;
   14805: out<=0;
   14806: out<=0;
   14807: out<=1;
   14808: out<=0;
   14809: out<=1;
   14810: out<=0;
   14811: out<=1;
   14812: out<=0;
   14813: out<=0;
   14814: out<=1;
   14815: out<=1;
   14816: out<=0;
   14817: out<=0;
   14818: out<=0;
   14819: out<=0;
   14820: out<=0;
   14821: out<=1;
   14822: out<=1;
   14823: out<=0;
   14824: out<=1;
   14825: out<=0;
   14826: out<=1;
   14827: out<=0;
   14828: out<=1;
   14829: out<=1;
   14830: out<=0;
   14831: out<=0;
   14832: out<=0;
   14833: out<=0;
   14834: out<=0;
   14835: out<=0;
   14836: out<=0;
   14837: out<=1;
   14838: out<=1;
   14839: out<=0;
   14840: out<=1;
   14841: out<=0;
   14842: out<=1;
   14843: out<=0;
   14844: out<=1;
   14845: out<=1;
   14846: out<=0;
   14847: out<=0;
   14848: out<=0;
   14849: out<=0;
   14850: out<=1;
   14851: out<=1;
   14852: out<=0;
   14853: out<=1;
   14854: out<=0;
   14855: out<=1;
   14856: out<=0;
   14857: out<=1;
   14858: out<=1;
   14859: out<=0;
   14860: out<=0;
   14861: out<=0;
   14862: out<=0;
   14863: out<=0;
   14864: out<=0;
   14865: out<=0;
   14866: out<=1;
   14867: out<=1;
   14868: out<=0;
   14869: out<=1;
   14870: out<=0;
   14871: out<=1;
   14872: out<=0;
   14873: out<=1;
   14874: out<=1;
   14875: out<=0;
   14876: out<=0;
   14877: out<=0;
   14878: out<=0;
   14879: out<=0;
   14880: out<=1;
   14881: out<=1;
   14882: out<=0;
   14883: out<=0;
   14884: out<=1;
   14885: out<=0;
   14886: out<=1;
   14887: out<=0;
   14888: out<=1;
   14889: out<=0;
   14890: out<=0;
   14891: out<=1;
   14892: out<=1;
   14893: out<=1;
   14894: out<=1;
   14895: out<=1;
   14896: out<=1;
   14897: out<=1;
   14898: out<=0;
   14899: out<=0;
   14900: out<=1;
   14901: out<=0;
   14902: out<=1;
   14903: out<=0;
   14904: out<=1;
   14905: out<=0;
   14906: out<=0;
   14907: out<=1;
   14908: out<=1;
   14909: out<=1;
   14910: out<=1;
   14911: out<=1;
   14912: out<=1;
   14913: out<=1;
   14914: out<=0;
   14915: out<=0;
   14916: out<=1;
   14917: out<=0;
   14918: out<=1;
   14919: out<=0;
   14920: out<=1;
   14921: out<=0;
   14922: out<=0;
   14923: out<=1;
   14924: out<=1;
   14925: out<=1;
   14926: out<=1;
   14927: out<=1;
   14928: out<=0;
   14929: out<=0;
   14930: out<=1;
   14931: out<=1;
   14932: out<=0;
   14933: out<=1;
   14934: out<=0;
   14935: out<=1;
   14936: out<=0;
   14937: out<=1;
   14938: out<=1;
   14939: out<=0;
   14940: out<=0;
   14941: out<=0;
   14942: out<=0;
   14943: out<=0;
   14944: out<=1;
   14945: out<=1;
   14946: out<=0;
   14947: out<=0;
   14948: out<=1;
   14949: out<=0;
   14950: out<=1;
   14951: out<=0;
   14952: out<=1;
   14953: out<=0;
   14954: out<=0;
   14955: out<=1;
   14956: out<=1;
   14957: out<=1;
   14958: out<=1;
   14959: out<=1;
   14960: out<=0;
   14961: out<=0;
   14962: out<=1;
   14963: out<=1;
   14964: out<=0;
   14965: out<=1;
   14966: out<=0;
   14967: out<=1;
   14968: out<=0;
   14969: out<=1;
   14970: out<=1;
   14971: out<=0;
   14972: out<=0;
   14973: out<=0;
   14974: out<=0;
   14975: out<=0;
   14976: out<=1;
   14977: out<=1;
   14978: out<=0;
   14979: out<=0;
   14980: out<=1;
   14981: out<=0;
   14982: out<=1;
   14983: out<=0;
   14984: out<=1;
   14985: out<=0;
   14986: out<=0;
   14987: out<=1;
   14988: out<=1;
   14989: out<=1;
   14990: out<=1;
   14991: out<=1;
   14992: out<=0;
   14993: out<=0;
   14994: out<=1;
   14995: out<=1;
   14996: out<=0;
   14997: out<=1;
   14998: out<=0;
   14999: out<=1;
   15000: out<=0;
   15001: out<=1;
   15002: out<=1;
   15003: out<=0;
   15004: out<=0;
   15005: out<=0;
   15006: out<=0;
   15007: out<=0;
   15008: out<=0;
   15009: out<=0;
   15010: out<=1;
   15011: out<=1;
   15012: out<=0;
   15013: out<=1;
   15014: out<=0;
   15015: out<=1;
   15016: out<=0;
   15017: out<=1;
   15018: out<=1;
   15019: out<=0;
   15020: out<=0;
   15021: out<=0;
   15022: out<=0;
   15023: out<=0;
   15024: out<=1;
   15025: out<=1;
   15026: out<=0;
   15027: out<=0;
   15028: out<=1;
   15029: out<=0;
   15030: out<=1;
   15031: out<=0;
   15032: out<=1;
   15033: out<=0;
   15034: out<=0;
   15035: out<=1;
   15036: out<=1;
   15037: out<=1;
   15038: out<=1;
   15039: out<=1;
   15040: out<=0;
   15041: out<=0;
   15042: out<=1;
   15043: out<=1;
   15044: out<=0;
   15045: out<=1;
   15046: out<=0;
   15047: out<=1;
   15048: out<=0;
   15049: out<=1;
   15050: out<=1;
   15051: out<=0;
   15052: out<=0;
   15053: out<=0;
   15054: out<=0;
   15055: out<=0;
   15056: out<=0;
   15057: out<=0;
   15058: out<=1;
   15059: out<=1;
   15060: out<=0;
   15061: out<=1;
   15062: out<=0;
   15063: out<=1;
   15064: out<=0;
   15065: out<=1;
   15066: out<=1;
   15067: out<=0;
   15068: out<=0;
   15069: out<=0;
   15070: out<=0;
   15071: out<=0;
   15072: out<=0;
   15073: out<=0;
   15074: out<=1;
   15075: out<=1;
   15076: out<=0;
   15077: out<=1;
   15078: out<=0;
   15079: out<=1;
   15080: out<=0;
   15081: out<=1;
   15082: out<=1;
   15083: out<=0;
   15084: out<=0;
   15085: out<=0;
   15086: out<=0;
   15087: out<=0;
   15088: out<=0;
   15089: out<=0;
   15090: out<=1;
   15091: out<=1;
   15092: out<=0;
   15093: out<=1;
   15094: out<=0;
   15095: out<=1;
   15096: out<=0;
   15097: out<=1;
   15098: out<=1;
   15099: out<=0;
   15100: out<=0;
   15101: out<=0;
   15102: out<=0;
   15103: out<=0;
   15104: out<=1;
   15105: out<=0;
   15106: out<=1;
   15107: out<=0;
   15108: out<=0;
   15109: out<=0;
   15110: out<=1;
   15111: out<=1;
   15112: out<=0;
   15113: out<=0;
   15114: out<=0;
   15115: out<=0;
   15116: out<=1;
   15117: out<=0;
   15118: out<=0;
   15119: out<=1;
   15120: out<=0;
   15121: out<=1;
   15122: out<=0;
   15123: out<=1;
   15124: out<=1;
   15125: out<=1;
   15126: out<=0;
   15127: out<=0;
   15128: out<=1;
   15129: out<=1;
   15130: out<=1;
   15131: out<=1;
   15132: out<=0;
   15133: out<=1;
   15134: out<=1;
   15135: out<=0;
   15136: out<=1;
   15137: out<=0;
   15138: out<=1;
   15139: out<=0;
   15140: out<=0;
   15141: out<=0;
   15142: out<=1;
   15143: out<=1;
   15144: out<=0;
   15145: out<=0;
   15146: out<=0;
   15147: out<=0;
   15148: out<=1;
   15149: out<=0;
   15150: out<=0;
   15151: out<=1;
   15152: out<=0;
   15153: out<=1;
   15154: out<=0;
   15155: out<=1;
   15156: out<=1;
   15157: out<=1;
   15158: out<=0;
   15159: out<=0;
   15160: out<=1;
   15161: out<=1;
   15162: out<=1;
   15163: out<=1;
   15164: out<=0;
   15165: out<=1;
   15166: out<=1;
   15167: out<=0;
   15168: out<=0;
   15169: out<=1;
   15170: out<=0;
   15171: out<=1;
   15172: out<=1;
   15173: out<=1;
   15174: out<=0;
   15175: out<=0;
   15176: out<=1;
   15177: out<=1;
   15178: out<=1;
   15179: out<=1;
   15180: out<=0;
   15181: out<=1;
   15182: out<=1;
   15183: out<=0;
   15184: out<=0;
   15185: out<=1;
   15186: out<=0;
   15187: out<=1;
   15188: out<=1;
   15189: out<=1;
   15190: out<=0;
   15191: out<=0;
   15192: out<=1;
   15193: out<=1;
   15194: out<=1;
   15195: out<=1;
   15196: out<=0;
   15197: out<=1;
   15198: out<=1;
   15199: out<=0;
   15200: out<=1;
   15201: out<=0;
   15202: out<=1;
   15203: out<=0;
   15204: out<=0;
   15205: out<=0;
   15206: out<=1;
   15207: out<=1;
   15208: out<=0;
   15209: out<=0;
   15210: out<=0;
   15211: out<=0;
   15212: out<=1;
   15213: out<=0;
   15214: out<=0;
   15215: out<=1;
   15216: out<=1;
   15217: out<=0;
   15218: out<=1;
   15219: out<=0;
   15220: out<=0;
   15221: out<=0;
   15222: out<=1;
   15223: out<=1;
   15224: out<=0;
   15225: out<=0;
   15226: out<=0;
   15227: out<=0;
   15228: out<=1;
   15229: out<=0;
   15230: out<=0;
   15231: out<=1;
   15232: out<=0;
   15233: out<=1;
   15234: out<=0;
   15235: out<=1;
   15236: out<=1;
   15237: out<=1;
   15238: out<=0;
   15239: out<=0;
   15240: out<=1;
   15241: out<=1;
   15242: out<=1;
   15243: out<=1;
   15244: out<=0;
   15245: out<=1;
   15246: out<=1;
   15247: out<=0;
   15248: out<=0;
   15249: out<=1;
   15250: out<=0;
   15251: out<=1;
   15252: out<=1;
   15253: out<=1;
   15254: out<=0;
   15255: out<=0;
   15256: out<=1;
   15257: out<=1;
   15258: out<=1;
   15259: out<=1;
   15260: out<=0;
   15261: out<=1;
   15262: out<=1;
   15263: out<=0;
   15264: out<=0;
   15265: out<=1;
   15266: out<=0;
   15267: out<=1;
   15268: out<=1;
   15269: out<=1;
   15270: out<=0;
   15271: out<=0;
   15272: out<=1;
   15273: out<=1;
   15274: out<=1;
   15275: out<=1;
   15276: out<=0;
   15277: out<=1;
   15278: out<=1;
   15279: out<=0;
   15280: out<=0;
   15281: out<=1;
   15282: out<=0;
   15283: out<=1;
   15284: out<=1;
   15285: out<=1;
   15286: out<=0;
   15287: out<=0;
   15288: out<=1;
   15289: out<=1;
   15290: out<=1;
   15291: out<=1;
   15292: out<=0;
   15293: out<=1;
   15294: out<=1;
   15295: out<=0;
   15296: out<=1;
   15297: out<=0;
   15298: out<=1;
   15299: out<=0;
   15300: out<=0;
   15301: out<=0;
   15302: out<=1;
   15303: out<=1;
   15304: out<=0;
   15305: out<=0;
   15306: out<=0;
   15307: out<=0;
   15308: out<=1;
   15309: out<=0;
   15310: out<=0;
   15311: out<=1;
   15312: out<=0;
   15313: out<=1;
   15314: out<=0;
   15315: out<=1;
   15316: out<=1;
   15317: out<=1;
   15318: out<=0;
   15319: out<=0;
   15320: out<=1;
   15321: out<=1;
   15322: out<=1;
   15323: out<=1;
   15324: out<=0;
   15325: out<=1;
   15326: out<=1;
   15327: out<=0;
   15328: out<=0;
   15329: out<=1;
   15330: out<=0;
   15331: out<=1;
   15332: out<=1;
   15333: out<=1;
   15334: out<=0;
   15335: out<=0;
   15336: out<=1;
   15337: out<=1;
   15338: out<=1;
   15339: out<=1;
   15340: out<=0;
   15341: out<=1;
   15342: out<=1;
   15343: out<=0;
   15344: out<=1;
   15345: out<=0;
   15346: out<=1;
   15347: out<=0;
   15348: out<=0;
   15349: out<=0;
   15350: out<=1;
   15351: out<=1;
   15352: out<=0;
   15353: out<=0;
   15354: out<=0;
   15355: out<=0;
   15356: out<=1;
   15357: out<=0;
   15358: out<=0;
   15359: out<=1;
   15360: out<=0;
   15361: out<=0;
   15362: out<=0;
   15363: out<=0;
   15364: out<=1;
   15365: out<=0;
   15366: out<=0;
   15367: out<=1;
   15368: out<=0;
   15369: out<=1;
   15370: out<=0;
   15371: out<=1;
   15372: out<=1;
   15373: out<=1;
   15374: out<=0;
   15375: out<=0;
   15376: out<=1;
   15377: out<=1;
   15378: out<=1;
   15379: out<=1;
   15380: out<=0;
   15381: out<=1;
   15382: out<=1;
   15383: out<=0;
   15384: out<=1;
   15385: out<=0;
   15386: out<=1;
   15387: out<=0;
   15388: out<=0;
   15389: out<=0;
   15390: out<=1;
   15391: out<=1;
   15392: out<=1;
   15393: out<=1;
   15394: out<=1;
   15395: out<=1;
   15396: out<=0;
   15397: out<=1;
   15398: out<=1;
   15399: out<=0;
   15400: out<=1;
   15401: out<=0;
   15402: out<=1;
   15403: out<=0;
   15404: out<=0;
   15405: out<=0;
   15406: out<=1;
   15407: out<=1;
   15408: out<=0;
   15409: out<=0;
   15410: out<=0;
   15411: out<=0;
   15412: out<=1;
   15413: out<=0;
   15414: out<=0;
   15415: out<=1;
   15416: out<=0;
   15417: out<=1;
   15418: out<=0;
   15419: out<=1;
   15420: out<=1;
   15421: out<=1;
   15422: out<=0;
   15423: out<=0;
   15424: out<=1;
   15425: out<=1;
   15426: out<=1;
   15427: out<=1;
   15428: out<=0;
   15429: out<=1;
   15430: out<=1;
   15431: out<=0;
   15432: out<=1;
   15433: out<=0;
   15434: out<=1;
   15435: out<=0;
   15436: out<=0;
   15437: out<=0;
   15438: out<=1;
   15439: out<=1;
   15440: out<=1;
   15441: out<=1;
   15442: out<=1;
   15443: out<=1;
   15444: out<=0;
   15445: out<=1;
   15446: out<=1;
   15447: out<=0;
   15448: out<=1;
   15449: out<=0;
   15450: out<=1;
   15451: out<=0;
   15452: out<=0;
   15453: out<=0;
   15454: out<=1;
   15455: out<=1;
   15456: out<=1;
   15457: out<=1;
   15458: out<=1;
   15459: out<=1;
   15460: out<=0;
   15461: out<=1;
   15462: out<=1;
   15463: out<=0;
   15464: out<=1;
   15465: out<=0;
   15466: out<=1;
   15467: out<=0;
   15468: out<=0;
   15469: out<=0;
   15470: out<=1;
   15471: out<=1;
   15472: out<=1;
   15473: out<=1;
   15474: out<=1;
   15475: out<=1;
   15476: out<=0;
   15477: out<=1;
   15478: out<=1;
   15479: out<=0;
   15480: out<=1;
   15481: out<=0;
   15482: out<=1;
   15483: out<=0;
   15484: out<=0;
   15485: out<=0;
   15486: out<=1;
   15487: out<=1;
   15488: out<=1;
   15489: out<=1;
   15490: out<=1;
   15491: out<=1;
   15492: out<=0;
   15493: out<=1;
   15494: out<=1;
   15495: out<=0;
   15496: out<=1;
   15497: out<=0;
   15498: out<=1;
   15499: out<=0;
   15500: out<=0;
   15501: out<=0;
   15502: out<=1;
   15503: out<=1;
   15504: out<=1;
   15505: out<=1;
   15506: out<=1;
   15507: out<=1;
   15508: out<=0;
   15509: out<=1;
   15510: out<=1;
   15511: out<=0;
   15512: out<=1;
   15513: out<=0;
   15514: out<=1;
   15515: out<=0;
   15516: out<=0;
   15517: out<=0;
   15518: out<=1;
   15519: out<=1;
   15520: out<=0;
   15521: out<=0;
   15522: out<=0;
   15523: out<=0;
   15524: out<=1;
   15525: out<=0;
   15526: out<=0;
   15527: out<=1;
   15528: out<=0;
   15529: out<=1;
   15530: out<=0;
   15531: out<=1;
   15532: out<=1;
   15533: out<=1;
   15534: out<=0;
   15535: out<=0;
   15536: out<=0;
   15537: out<=0;
   15538: out<=0;
   15539: out<=0;
   15540: out<=1;
   15541: out<=0;
   15542: out<=0;
   15543: out<=1;
   15544: out<=0;
   15545: out<=1;
   15546: out<=0;
   15547: out<=1;
   15548: out<=1;
   15549: out<=1;
   15550: out<=0;
   15551: out<=0;
   15552: out<=0;
   15553: out<=0;
   15554: out<=0;
   15555: out<=0;
   15556: out<=1;
   15557: out<=0;
   15558: out<=0;
   15559: out<=1;
   15560: out<=0;
   15561: out<=1;
   15562: out<=0;
   15563: out<=1;
   15564: out<=1;
   15565: out<=1;
   15566: out<=0;
   15567: out<=0;
   15568: out<=1;
   15569: out<=1;
   15570: out<=1;
   15571: out<=1;
   15572: out<=0;
   15573: out<=1;
   15574: out<=1;
   15575: out<=0;
   15576: out<=1;
   15577: out<=0;
   15578: out<=1;
   15579: out<=0;
   15580: out<=0;
   15581: out<=0;
   15582: out<=1;
   15583: out<=1;
   15584: out<=0;
   15585: out<=0;
   15586: out<=0;
   15587: out<=0;
   15588: out<=1;
   15589: out<=0;
   15590: out<=0;
   15591: out<=1;
   15592: out<=0;
   15593: out<=1;
   15594: out<=0;
   15595: out<=1;
   15596: out<=1;
   15597: out<=1;
   15598: out<=0;
   15599: out<=0;
   15600: out<=1;
   15601: out<=1;
   15602: out<=1;
   15603: out<=1;
   15604: out<=0;
   15605: out<=1;
   15606: out<=1;
   15607: out<=0;
   15608: out<=1;
   15609: out<=0;
   15610: out<=1;
   15611: out<=0;
   15612: out<=0;
   15613: out<=0;
   15614: out<=1;
   15615: out<=1;
   15616: out<=0;
   15617: out<=1;
   15618: out<=1;
   15619: out<=0;
   15620: out<=0;
   15621: out<=0;
   15622: out<=0;
   15623: out<=0;
   15624: out<=1;
   15625: out<=1;
   15626: out<=0;
   15627: out<=0;
   15628: out<=1;
   15629: out<=0;
   15630: out<=1;
   15631: out<=0;
   15632: out<=0;
   15633: out<=1;
   15634: out<=1;
   15635: out<=0;
   15636: out<=0;
   15637: out<=0;
   15638: out<=0;
   15639: out<=0;
   15640: out<=1;
   15641: out<=1;
   15642: out<=0;
   15643: out<=0;
   15644: out<=1;
   15645: out<=0;
   15646: out<=1;
   15647: out<=0;
   15648: out<=0;
   15649: out<=1;
   15650: out<=1;
   15651: out<=0;
   15652: out<=0;
   15653: out<=0;
   15654: out<=0;
   15655: out<=0;
   15656: out<=1;
   15657: out<=1;
   15658: out<=0;
   15659: out<=0;
   15660: out<=1;
   15661: out<=0;
   15662: out<=1;
   15663: out<=0;
   15664: out<=0;
   15665: out<=1;
   15666: out<=1;
   15667: out<=0;
   15668: out<=0;
   15669: out<=0;
   15670: out<=0;
   15671: out<=0;
   15672: out<=1;
   15673: out<=1;
   15674: out<=0;
   15675: out<=0;
   15676: out<=1;
   15677: out<=0;
   15678: out<=1;
   15679: out<=0;
   15680: out<=1;
   15681: out<=0;
   15682: out<=0;
   15683: out<=1;
   15684: out<=1;
   15685: out<=1;
   15686: out<=1;
   15687: out<=1;
   15688: out<=0;
   15689: out<=0;
   15690: out<=1;
   15691: out<=1;
   15692: out<=0;
   15693: out<=1;
   15694: out<=0;
   15695: out<=1;
   15696: out<=0;
   15697: out<=1;
   15698: out<=1;
   15699: out<=0;
   15700: out<=0;
   15701: out<=0;
   15702: out<=0;
   15703: out<=0;
   15704: out<=1;
   15705: out<=1;
   15706: out<=0;
   15707: out<=0;
   15708: out<=1;
   15709: out<=0;
   15710: out<=1;
   15711: out<=0;
   15712: out<=0;
   15713: out<=1;
   15714: out<=1;
   15715: out<=0;
   15716: out<=0;
   15717: out<=0;
   15718: out<=0;
   15719: out<=0;
   15720: out<=1;
   15721: out<=1;
   15722: out<=0;
   15723: out<=0;
   15724: out<=1;
   15725: out<=0;
   15726: out<=1;
   15727: out<=0;
   15728: out<=1;
   15729: out<=0;
   15730: out<=0;
   15731: out<=1;
   15732: out<=1;
   15733: out<=1;
   15734: out<=1;
   15735: out<=1;
   15736: out<=0;
   15737: out<=0;
   15738: out<=1;
   15739: out<=1;
   15740: out<=0;
   15741: out<=1;
   15742: out<=0;
   15743: out<=1;
   15744: out<=1;
   15745: out<=0;
   15746: out<=0;
   15747: out<=1;
   15748: out<=1;
   15749: out<=1;
   15750: out<=1;
   15751: out<=1;
   15752: out<=0;
   15753: out<=0;
   15754: out<=1;
   15755: out<=1;
   15756: out<=0;
   15757: out<=1;
   15758: out<=0;
   15759: out<=1;
   15760: out<=0;
   15761: out<=1;
   15762: out<=1;
   15763: out<=0;
   15764: out<=0;
   15765: out<=0;
   15766: out<=0;
   15767: out<=0;
   15768: out<=1;
   15769: out<=1;
   15770: out<=0;
   15771: out<=0;
   15772: out<=1;
   15773: out<=0;
   15774: out<=1;
   15775: out<=0;
   15776: out<=1;
   15777: out<=0;
   15778: out<=0;
   15779: out<=1;
   15780: out<=1;
   15781: out<=1;
   15782: out<=1;
   15783: out<=1;
   15784: out<=0;
   15785: out<=0;
   15786: out<=1;
   15787: out<=1;
   15788: out<=0;
   15789: out<=1;
   15790: out<=0;
   15791: out<=1;
   15792: out<=0;
   15793: out<=1;
   15794: out<=1;
   15795: out<=0;
   15796: out<=0;
   15797: out<=0;
   15798: out<=0;
   15799: out<=0;
   15800: out<=1;
   15801: out<=1;
   15802: out<=0;
   15803: out<=0;
   15804: out<=1;
   15805: out<=0;
   15806: out<=1;
   15807: out<=0;
   15808: out<=0;
   15809: out<=1;
   15810: out<=1;
   15811: out<=0;
   15812: out<=0;
   15813: out<=0;
   15814: out<=0;
   15815: out<=0;
   15816: out<=1;
   15817: out<=1;
   15818: out<=0;
   15819: out<=0;
   15820: out<=1;
   15821: out<=0;
   15822: out<=1;
   15823: out<=0;
   15824: out<=0;
   15825: out<=1;
   15826: out<=1;
   15827: out<=0;
   15828: out<=0;
   15829: out<=0;
   15830: out<=0;
   15831: out<=0;
   15832: out<=1;
   15833: out<=1;
   15834: out<=0;
   15835: out<=0;
   15836: out<=1;
   15837: out<=0;
   15838: out<=1;
   15839: out<=0;
   15840: out<=1;
   15841: out<=0;
   15842: out<=0;
   15843: out<=1;
   15844: out<=1;
   15845: out<=1;
   15846: out<=1;
   15847: out<=1;
   15848: out<=0;
   15849: out<=0;
   15850: out<=1;
   15851: out<=1;
   15852: out<=0;
   15853: out<=1;
   15854: out<=0;
   15855: out<=1;
   15856: out<=1;
   15857: out<=0;
   15858: out<=0;
   15859: out<=1;
   15860: out<=1;
   15861: out<=1;
   15862: out<=1;
   15863: out<=1;
   15864: out<=0;
   15865: out<=0;
   15866: out<=1;
   15867: out<=1;
   15868: out<=0;
   15869: out<=1;
   15870: out<=0;
   15871: out<=1;
   15872: out<=1;
   15873: out<=0;
   15874: out<=1;
   15875: out<=0;
   15876: out<=1;
   15877: out<=1;
   15878: out<=0;
   15879: out<=0;
   15880: out<=1;
   15881: out<=1;
   15882: out<=1;
   15883: out<=1;
   15884: out<=1;
   15885: out<=0;
   15886: out<=0;
   15887: out<=1;
   15888: out<=1;
   15889: out<=0;
   15890: out<=1;
   15891: out<=0;
   15892: out<=1;
   15893: out<=1;
   15894: out<=0;
   15895: out<=0;
   15896: out<=1;
   15897: out<=1;
   15898: out<=1;
   15899: out<=1;
   15900: out<=1;
   15901: out<=0;
   15902: out<=0;
   15903: out<=1;
   15904: out<=0;
   15905: out<=1;
   15906: out<=0;
   15907: out<=1;
   15908: out<=0;
   15909: out<=0;
   15910: out<=1;
   15911: out<=1;
   15912: out<=0;
   15913: out<=0;
   15914: out<=0;
   15915: out<=0;
   15916: out<=0;
   15917: out<=1;
   15918: out<=1;
   15919: out<=0;
   15920: out<=0;
   15921: out<=1;
   15922: out<=0;
   15923: out<=1;
   15924: out<=0;
   15925: out<=0;
   15926: out<=1;
   15927: out<=1;
   15928: out<=0;
   15929: out<=0;
   15930: out<=0;
   15931: out<=0;
   15932: out<=0;
   15933: out<=1;
   15934: out<=1;
   15935: out<=0;
   15936: out<=0;
   15937: out<=1;
   15938: out<=0;
   15939: out<=1;
   15940: out<=0;
   15941: out<=0;
   15942: out<=1;
   15943: out<=1;
   15944: out<=0;
   15945: out<=0;
   15946: out<=0;
   15947: out<=0;
   15948: out<=0;
   15949: out<=1;
   15950: out<=1;
   15951: out<=0;
   15952: out<=1;
   15953: out<=0;
   15954: out<=1;
   15955: out<=0;
   15956: out<=1;
   15957: out<=1;
   15958: out<=0;
   15959: out<=0;
   15960: out<=1;
   15961: out<=1;
   15962: out<=1;
   15963: out<=1;
   15964: out<=1;
   15965: out<=0;
   15966: out<=0;
   15967: out<=1;
   15968: out<=0;
   15969: out<=1;
   15970: out<=0;
   15971: out<=1;
   15972: out<=0;
   15973: out<=0;
   15974: out<=1;
   15975: out<=1;
   15976: out<=0;
   15977: out<=0;
   15978: out<=0;
   15979: out<=0;
   15980: out<=0;
   15981: out<=1;
   15982: out<=1;
   15983: out<=0;
   15984: out<=1;
   15985: out<=0;
   15986: out<=1;
   15987: out<=0;
   15988: out<=1;
   15989: out<=1;
   15990: out<=0;
   15991: out<=0;
   15992: out<=1;
   15993: out<=1;
   15994: out<=1;
   15995: out<=1;
   15996: out<=1;
   15997: out<=0;
   15998: out<=0;
   15999: out<=1;
   16000: out<=0;
   16001: out<=1;
   16002: out<=0;
   16003: out<=1;
   16004: out<=0;
   16005: out<=0;
   16006: out<=1;
   16007: out<=1;
   16008: out<=0;
   16009: out<=0;
   16010: out<=0;
   16011: out<=0;
   16012: out<=0;
   16013: out<=1;
   16014: out<=1;
   16015: out<=0;
   16016: out<=1;
   16017: out<=0;
   16018: out<=1;
   16019: out<=0;
   16020: out<=1;
   16021: out<=1;
   16022: out<=0;
   16023: out<=0;
   16024: out<=1;
   16025: out<=1;
   16026: out<=1;
   16027: out<=1;
   16028: out<=1;
   16029: out<=0;
   16030: out<=0;
   16031: out<=1;
   16032: out<=1;
   16033: out<=0;
   16034: out<=1;
   16035: out<=0;
   16036: out<=1;
   16037: out<=1;
   16038: out<=0;
   16039: out<=0;
   16040: out<=1;
   16041: out<=1;
   16042: out<=1;
   16043: out<=1;
   16044: out<=1;
   16045: out<=0;
   16046: out<=0;
   16047: out<=1;
   16048: out<=0;
   16049: out<=1;
   16050: out<=0;
   16051: out<=1;
   16052: out<=0;
   16053: out<=0;
   16054: out<=1;
   16055: out<=1;
   16056: out<=0;
   16057: out<=0;
   16058: out<=0;
   16059: out<=0;
   16060: out<=0;
   16061: out<=1;
   16062: out<=1;
   16063: out<=0;
   16064: out<=1;
   16065: out<=0;
   16066: out<=1;
   16067: out<=0;
   16068: out<=1;
   16069: out<=1;
   16070: out<=0;
   16071: out<=0;
   16072: out<=1;
   16073: out<=1;
   16074: out<=1;
   16075: out<=1;
   16076: out<=1;
   16077: out<=0;
   16078: out<=0;
   16079: out<=1;
   16080: out<=1;
   16081: out<=0;
   16082: out<=1;
   16083: out<=0;
   16084: out<=1;
   16085: out<=1;
   16086: out<=0;
   16087: out<=0;
   16088: out<=1;
   16089: out<=1;
   16090: out<=1;
   16091: out<=1;
   16092: out<=1;
   16093: out<=0;
   16094: out<=0;
   16095: out<=1;
   16096: out<=1;
   16097: out<=0;
   16098: out<=1;
   16099: out<=0;
   16100: out<=1;
   16101: out<=1;
   16102: out<=0;
   16103: out<=0;
   16104: out<=1;
   16105: out<=1;
   16106: out<=1;
   16107: out<=1;
   16108: out<=1;
   16109: out<=0;
   16110: out<=0;
   16111: out<=1;
   16112: out<=1;
   16113: out<=0;
   16114: out<=1;
   16115: out<=0;
   16116: out<=1;
   16117: out<=1;
   16118: out<=0;
   16119: out<=0;
   16120: out<=1;
   16121: out<=1;
   16122: out<=1;
   16123: out<=1;
   16124: out<=1;
   16125: out<=0;
   16126: out<=0;
   16127: out<=1;
   16128: out<=1;
   16129: out<=1;
   16130: out<=0;
   16131: out<=0;
   16132: out<=0;
   16133: out<=1;
   16134: out<=0;
   16135: out<=1;
   16136: out<=0;
   16137: out<=1;
   16138: out<=1;
   16139: out<=0;
   16140: out<=1;
   16141: out<=1;
   16142: out<=1;
   16143: out<=1;
   16144: out<=0;
   16145: out<=0;
   16146: out<=1;
   16147: out<=1;
   16148: out<=1;
   16149: out<=0;
   16150: out<=1;
   16151: out<=0;
   16152: out<=1;
   16153: out<=0;
   16154: out<=0;
   16155: out<=1;
   16156: out<=0;
   16157: out<=0;
   16158: out<=0;
   16159: out<=0;
   16160: out<=1;
   16161: out<=1;
   16162: out<=0;
   16163: out<=0;
   16164: out<=0;
   16165: out<=1;
   16166: out<=0;
   16167: out<=1;
   16168: out<=0;
   16169: out<=1;
   16170: out<=1;
   16171: out<=0;
   16172: out<=1;
   16173: out<=1;
   16174: out<=1;
   16175: out<=1;
   16176: out<=0;
   16177: out<=0;
   16178: out<=1;
   16179: out<=1;
   16180: out<=1;
   16181: out<=0;
   16182: out<=1;
   16183: out<=0;
   16184: out<=1;
   16185: out<=0;
   16186: out<=0;
   16187: out<=1;
   16188: out<=0;
   16189: out<=0;
   16190: out<=0;
   16191: out<=0;
   16192: out<=0;
   16193: out<=0;
   16194: out<=1;
   16195: out<=1;
   16196: out<=1;
   16197: out<=0;
   16198: out<=1;
   16199: out<=0;
   16200: out<=1;
   16201: out<=0;
   16202: out<=0;
   16203: out<=1;
   16204: out<=0;
   16205: out<=0;
   16206: out<=0;
   16207: out<=0;
   16208: out<=0;
   16209: out<=0;
   16210: out<=1;
   16211: out<=1;
   16212: out<=1;
   16213: out<=0;
   16214: out<=1;
   16215: out<=0;
   16216: out<=1;
   16217: out<=0;
   16218: out<=0;
   16219: out<=1;
   16220: out<=0;
   16221: out<=0;
   16222: out<=0;
   16223: out<=0;
   16224: out<=1;
   16225: out<=1;
   16226: out<=0;
   16227: out<=0;
   16228: out<=0;
   16229: out<=1;
   16230: out<=0;
   16231: out<=1;
   16232: out<=0;
   16233: out<=1;
   16234: out<=1;
   16235: out<=0;
   16236: out<=1;
   16237: out<=1;
   16238: out<=1;
   16239: out<=1;
   16240: out<=1;
   16241: out<=1;
   16242: out<=0;
   16243: out<=0;
   16244: out<=0;
   16245: out<=1;
   16246: out<=0;
   16247: out<=1;
   16248: out<=0;
   16249: out<=1;
   16250: out<=1;
   16251: out<=0;
   16252: out<=1;
   16253: out<=1;
   16254: out<=1;
   16255: out<=1;
   16256: out<=0;
   16257: out<=0;
   16258: out<=1;
   16259: out<=1;
   16260: out<=1;
   16261: out<=0;
   16262: out<=1;
   16263: out<=0;
   16264: out<=1;
   16265: out<=0;
   16266: out<=0;
   16267: out<=1;
   16268: out<=0;
   16269: out<=0;
   16270: out<=0;
   16271: out<=0;
   16272: out<=0;
   16273: out<=0;
   16274: out<=1;
   16275: out<=1;
   16276: out<=1;
   16277: out<=0;
   16278: out<=1;
   16279: out<=0;
   16280: out<=1;
   16281: out<=0;
   16282: out<=0;
   16283: out<=1;
   16284: out<=0;
   16285: out<=0;
   16286: out<=0;
   16287: out<=0;
   16288: out<=0;
   16289: out<=0;
   16290: out<=1;
   16291: out<=1;
   16292: out<=1;
   16293: out<=0;
   16294: out<=1;
   16295: out<=0;
   16296: out<=1;
   16297: out<=0;
   16298: out<=0;
   16299: out<=1;
   16300: out<=0;
   16301: out<=0;
   16302: out<=0;
   16303: out<=0;
   16304: out<=0;
   16305: out<=0;
   16306: out<=1;
   16307: out<=1;
   16308: out<=1;
   16309: out<=0;
   16310: out<=1;
   16311: out<=0;
   16312: out<=1;
   16313: out<=0;
   16314: out<=0;
   16315: out<=1;
   16316: out<=0;
   16317: out<=0;
   16318: out<=0;
   16319: out<=0;
   16320: out<=1;
   16321: out<=1;
   16322: out<=0;
   16323: out<=0;
   16324: out<=0;
   16325: out<=1;
   16326: out<=0;
   16327: out<=1;
   16328: out<=0;
   16329: out<=1;
   16330: out<=1;
   16331: out<=0;
   16332: out<=1;
   16333: out<=1;
   16334: out<=1;
   16335: out<=1;
   16336: out<=0;
   16337: out<=0;
   16338: out<=1;
   16339: out<=1;
   16340: out<=1;
   16341: out<=0;
   16342: out<=1;
   16343: out<=0;
   16344: out<=1;
   16345: out<=0;
   16346: out<=0;
   16347: out<=1;
   16348: out<=0;
   16349: out<=0;
   16350: out<=0;
   16351: out<=0;
   16352: out<=0;
   16353: out<=0;
   16354: out<=1;
   16355: out<=1;
   16356: out<=1;
   16357: out<=0;
   16358: out<=1;
   16359: out<=0;
   16360: out<=1;
   16361: out<=0;
   16362: out<=0;
   16363: out<=1;
   16364: out<=0;
   16365: out<=0;
   16366: out<=0;
   16367: out<=0;
   16368: out<=1;
   16369: out<=1;
   16370: out<=0;
   16371: out<=0;
   16372: out<=0;
   16373: out<=1;
   16374: out<=0;
   16375: out<=1;
   16376: out<=0;
   16377: out<=1;
   16378: out<=1;
   16379: out<=0;
   16380: out<=1;
   16381: out<=1;
   16382: out<=1;
   16383: out<=1;
   16384: out<=0;
   16385: out<=0;
   16386: out<=0;
   16387: out<=0;
   16388: out<=1;
   16389: out<=0;
   16390: out<=0;
   16391: out<=1;
   16392: out<=0;
   16393: out<=1;
   16394: out<=0;
   16395: out<=1;
   16396: out<=1;
   16397: out<=1;
   16398: out<=0;
   16399: out<=0;
   16400: out<=0;
   16401: out<=0;
   16402: out<=0;
   16403: out<=0;
   16404: out<=1;
   16405: out<=0;
   16406: out<=0;
   16407: out<=1;
   16408: out<=0;
   16409: out<=1;
   16410: out<=0;
   16411: out<=1;
   16412: out<=1;
   16413: out<=1;
   16414: out<=0;
   16415: out<=0;
   16416: out<=1;
   16417: out<=1;
   16418: out<=1;
   16419: out<=1;
   16420: out<=0;
   16421: out<=1;
   16422: out<=1;
   16423: out<=0;
   16424: out<=1;
   16425: out<=0;
   16426: out<=1;
   16427: out<=0;
   16428: out<=0;
   16429: out<=0;
   16430: out<=1;
   16431: out<=1;
   16432: out<=1;
   16433: out<=1;
   16434: out<=1;
   16435: out<=1;
   16436: out<=0;
   16437: out<=1;
   16438: out<=1;
   16439: out<=0;
   16440: out<=1;
   16441: out<=0;
   16442: out<=1;
   16443: out<=0;
   16444: out<=0;
   16445: out<=0;
   16446: out<=1;
   16447: out<=1;
   16448: out<=1;
   16449: out<=1;
   16450: out<=1;
   16451: out<=1;
   16452: out<=0;
   16453: out<=1;
   16454: out<=1;
   16455: out<=0;
   16456: out<=1;
   16457: out<=0;
   16458: out<=1;
   16459: out<=0;
   16460: out<=0;
   16461: out<=0;
   16462: out<=1;
   16463: out<=1;
   16464: out<=0;
   16465: out<=0;
   16466: out<=0;
   16467: out<=0;
   16468: out<=1;
   16469: out<=0;
   16470: out<=0;
   16471: out<=1;
   16472: out<=0;
   16473: out<=1;
   16474: out<=0;
   16475: out<=1;
   16476: out<=1;
   16477: out<=1;
   16478: out<=0;
   16479: out<=0;
   16480: out<=1;
   16481: out<=1;
   16482: out<=1;
   16483: out<=1;
   16484: out<=0;
   16485: out<=1;
   16486: out<=1;
   16487: out<=0;
   16488: out<=1;
   16489: out<=0;
   16490: out<=1;
   16491: out<=0;
   16492: out<=0;
   16493: out<=0;
   16494: out<=1;
   16495: out<=1;
   16496: out<=0;
   16497: out<=0;
   16498: out<=0;
   16499: out<=0;
   16500: out<=1;
   16501: out<=0;
   16502: out<=0;
   16503: out<=1;
   16504: out<=0;
   16505: out<=1;
   16506: out<=0;
   16507: out<=1;
   16508: out<=1;
   16509: out<=1;
   16510: out<=0;
   16511: out<=0;
   16512: out<=0;
   16513: out<=0;
   16514: out<=0;
   16515: out<=0;
   16516: out<=1;
   16517: out<=0;
   16518: out<=0;
   16519: out<=1;
   16520: out<=0;
   16521: out<=1;
   16522: out<=0;
   16523: out<=1;
   16524: out<=1;
   16525: out<=1;
   16526: out<=0;
   16527: out<=0;
   16528: out<=1;
   16529: out<=1;
   16530: out<=1;
   16531: out<=1;
   16532: out<=0;
   16533: out<=1;
   16534: out<=1;
   16535: out<=0;
   16536: out<=1;
   16537: out<=0;
   16538: out<=1;
   16539: out<=0;
   16540: out<=0;
   16541: out<=0;
   16542: out<=1;
   16543: out<=1;
   16544: out<=1;
   16545: out<=1;
   16546: out<=1;
   16547: out<=1;
   16548: out<=0;
   16549: out<=1;
   16550: out<=1;
   16551: out<=0;
   16552: out<=1;
   16553: out<=0;
   16554: out<=1;
   16555: out<=0;
   16556: out<=0;
   16557: out<=0;
   16558: out<=1;
   16559: out<=1;
   16560: out<=0;
   16561: out<=0;
   16562: out<=0;
   16563: out<=0;
   16564: out<=1;
   16565: out<=0;
   16566: out<=0;
   16567: out<=1;
   16568: out<=0;
   16569: out<=1;
   16570: out<=0;
   16571: out<=1;
   16572: out<=1;
   16573: out<=1;
   16574: out<=0;
   16575: out<=0;
   16576: out<=1;
   16577: out<=1;
   16578: out<=1;
   16579: out<=1;
   16580: out<=0;
   16581: out<=1;
   16582: out<=1;
   16583: out<=0;
   16584: out<=1;
   16585: out<=0;
   16586: out<=1;
   16587: out<=0;
   16588: out<=0;
   16589: out<=0;
   16590: out<=1;
   16591: out<=1;
   16592: out<=1;
   16593: out<=1;
   16594: out<=1;
   16595: out<=1;
   16596: out<=0;
   16597: out<=1;
   16598: out<=1;
   16599: out<=0;
   16600: out<=1;
   16601: out<=0;
   16602: out<=1;
   16603: out<=0;
   16604: out<=0;
   16605: out<=0;
   16606: out<=1;
   16607: out<=1;
   16608: out<=1;
   16609: out<=1;
   16610: out<=1;
   16611: out<=1;
   16612: out<=0;
   16613: out<=1;
   16614: out<=1;
   16615: out<=0;
   16616: out<=1;
   16617: out<=0;
   16618: out<=1;
   16619: out<=0;
   16620: out<=0;
   16621: out<=0;
   16622: out<=1;
   16623: out<=1;
   16624: out<=1;
   16625: out<=1;
   16626: out<=1;
   16627: out<=1;
   16628: out<=0;
   16629: out<=1;
   16630: out<=1;
   16631: out<=0;
   16632: out<=1;
   16633: out<=0;
   16634: out<=1;
   16635: out<=0;
   16636: out<=0;
   16637: out<=0;
   16638: out<=1;
   16639: out<=1;
   16640: out<=0;
   16641: out<=1;
   16642: out<=1;
   16643: out<=0;
   16644: out<=0;
   16645: out<=0;
   16646: out<=0;
   16647: out<=0;
   16648: out<=1;
   16649: out<=1;
   16650: out<=0;
   16651: out<=0;
   16652: out<=1;
   16653: out<=0;
   16654: out<=1;
   16655: out<=0;
   16656: out<=1;
   16657: out<=0;
   16658: out<=0;
   16659: out<=1;
   16660: out<=1;
   16661: out<=1;
   16662: out<=1;
   16663: out<=1;
   16664: out<=0;
   16665: out<=0;
   16666: out<=1;
   16667: out<=1;
   16668: out<=0;
   16669: out<=1;
   16670: out<=0;
   16671: out<=1;
   16672: out<=0;
   16673: out<=1;
   16674: out<=1;
   16675: out<=0;
   16676: out<=0;
   16677: out<=0;
   16678: out<=0;
   16679: out<=0;
   16680: out<=1;
   16681: out<=1;
   16682: out<=0;
   16683: out<=0;
   16684: out<=1;
   16685: out<=0;
   16686: out<=1;
   16687: out<=0;
   16688: out<=1;
   16689: out<=0;
   16690: out<=0;
   16691: out<=1;
   16692: out<=1;
   16693: out<=1;
   16694: out<=1;
   16695: out<=1;
   16696: out<=0;
   16697: out<=0;
   16698: out<=1;
   16699: out<=1;
   16700: out<=0;
   16701: out<=1;
   16702: out<=0;
   16703: out<=1;
   16704: out<=1;
   16705: out<=0;
   16706: out<=0;
   16707: out<=1;
   16708: out<=1;
   16709: out<=1;
   16710: out<=1;
   16711: out<=1;
   16712: out<=0;
   16713: out<=0;
   16714: out<=1;
   16715: out<=1;
   16716: out<=0;
   16717: out<=1;
   16718: out<=0;
   16719: out<=1;
   16720: out<=1;
   16721: out<=0;
   16722: out<=0;
   16723: out<=1;
   16724: out<=1;
   16725: out<=1;
   16726: out<=1;
   16727: out<=1;
   16728: out<=0;
   16729: out<=0;
   16730: out<=1;
   16731: out<=1;
   16732: out<=0;
   16733: out<=1;
   16734: out<=0;
   16735: out<=1;
   16736: out<=0;
   16737: out<=1;
   16738: out<=1;
   16739: out<=0;
   16740: out<=0;
   16741: out<=0;
   16742: out<=0;
   16743: out<=0;
   16744: out<=1;
   16745: out<=1;
   16746: out<=0;
   16747: out<=0;
   16748: out<=1;
   16749: out<=0;
   16750: out<=1;
   16751: out<=0;
   16752: out<=0;
   16753: out<=1;
   16754: out<=1;
   16755: out<=0;
   16756: out<=0;
   16757: out<=0;
   16758: out<=0;
   16759: out<=0;
   16760: out<=1;
   16761: out<=1;
   16762: out<=0;
   16763: out<=0;
   16764: out<=1;
   16765: out<=0;
   16766: out<=1;
   16767: out<=0;
   16768: out<=0;
   16769: out<=1;
   16770: out<=1;
   16771: out<=0;
   16772: out<=0;
   16773: out<=0;
   16774: out<=0;
   16775: out<=0;
   16776: out<=1;
   16777: out<=1;
   16778: out<=0;
   16779: out<=0;
   16780: out<=1;
   16781: out<=0;
   16782: out<=1;
   16783: out<=0;
   16784: out<=0;
   16785: out<=1;
   16786: out<=1;
   16787: out<=0;
   16788: out<=0;
   16789: out<=0;
   16790: out<=0;
   16791: out<=0;
   16792: out<=1;
   16793: out<=1;
   16794: out<=0;
   16795: out<=0;
   16796: out<=1;
   16797: out<=0;
   16798: out<=1;
   16799: out<=0;
   16800: out<=0;
   16801: out<=1;
   16802: out<=1;
   16803: out<=0;
   16804: out<=0;
   16805: out<=0;
   16806: out<=0;
   16807: out<=0;
   16808: out<=1;
   16809: out<=1;
   16810: out<=0;
   16811: out<=0;
   16812: out<=1;
   16813: out<=0;
   16814: out<=1;
   16815: out<=0;
   16816: out<=0;
   16817: out<=1;
   16818: out<=1;
   16819: out<=0;
   16820: out<=0;
   16821: out<=0;
   16822: out<=0;
   16823: out<=0;
   16824: out<=1;
   16825: out<=1;
   16826: out<=0;
   16827: out<=0;
   16828: out<=1;
   16829: out<=0;
   16830: out<=1;
   16831: out<=0;
   16832: out<=1;
   16833: out<=0;
   16834: out<=0;
   16835: out<=1;
   16836: out<=1;
   16837: out<=1;
   16838: out<=1;
   16839: out<=1;
   16840: out<=0;
   16841: out<=0;
   16842: out<=1;
   16843: out<=1;
   16844: out<=0;
   16845: out<=1;
   16846: out<=0;
   16847: out<=1;
   16848: out<=0;
   16849: out<=1;
   16850: out<=1;
   16851: out<=0;
   16852: out<=0;
   16853: out<=0;
   16854: out<=0;
   16855: out<=0;
   16856: out<=1;
   16857: out<=1;
   16858: out<=0;
   16859: out<=0;
   16860: out<=1;
   16861: out<=0;
   16862: out<=1;
   16863: out<=0;
   16864: out<=0;
   16865: out<=1;
   16866: out<=1;
   16867: out<=0;
   16868: out<=0;
   16869: out<=0;
   16870: out<=0;
   16871: out<=0;
   16872: out<=1;
   16873: out<=1;
   16874: out<=0;
   16875: out<=0;
   16876: out<=1;
   16877: out<=0;
   16878: out<=1;
   16879: out<=0;
   16880: out<=1;
   16881: out<=0;
   16882: out<=0;
   16883: out<=1;
   16884: out<=1;
   16885: out<=1;
   16886: out<=1;
   16887: out<=1;
   16888: out<=0;
   16889: out<=0;
   16890: out<=1;
   16891: out<=1;
   16892: out<=0;
   16893: out<=1;
   16894: out<=0;
   16895: out<=1;
   16896: out<=0;
   16897: out<=1;
   16898: out<=0;
   16899: out<=1;
   16900: out<=0;
   16901: out<=0;
   16902: out<=1;
   16903: out<=1;
   16904: out<=0;
   16905: out<=0;
   16906: out<=0;
   16907: out<=0;
   16908: out<=0;
   16909: out<=1;
   16910: out<=1;
   16911: out<=0;
   16912: out<=1;
   16913: out<=0;
   16914: out<=1;
   16915: out<=0;
   16916: out<=1;
   16917: out<=1;
   16918: out<=0;
   16919: out<=0;
   16920: out<=1;
   16921: out<=1;
   16922: out<=1;
   16923: out<=1;
   16924: out<=1;
   16925: out<=0;
   16926: out<=0;
   16927: out<=1;
   16928: out<=1;
   16929: out<=0;
   16930: out<=1;
   16931: out<=0;
   16932: out<=1;
   16933: out<=1;
   16934: out<=0;
   16935: out<=0;
   16936: out<=1;
   16937: out<=1;
   16938: out<=1;
   16939: out<=1;
   16940: out<=1;
   16941: out<=0;
   16942: out<=0;
   16943: out<=1;
   16944: out<=0;
   16945: out<=1;
   16946: out<=0;
   16947: out<=1;
   16948: out<=0;
   16949: out<=0;
   16950: out<=1;
   16951: out<=1;
   16952: out<=0;
   16953: out<=0;
   16954: out<=0;
   16955: out<=0;
   16956: out<=0;
   16957: out<=1;
   16958: out<=1;
   16959: out<=0;
   16960: out<=1;
   16961: out<=0;
   16962: out<=1;
   16963: out<=0;
   16964: out<=1;
   16965: out<=1;
   16966: out<=0;
   16967: out<=0;
   16968: out<=1;
   16969: out<=1;
   16970: out<=1;
   16971: out<=1;
   16972: out<=1;
   16973: out<=0;
   16974: out<=0;
   16975: out<=1;
   16976: out<=1;
   16977: out<=0;
   16978: out<=1;
   16979: out<=0;
   16980: out<=1;
   16981: out<=1;
   16982: out<=0;
   16983: out<=0;
   16984: out<=1;
   16985: out<=1;
   16986: out<=1;
   16987: out<=1;
   16988: out<=1;
   16989: out<=0;
   16990: out<=0;
   16991: out<=1;
   16992: out<=1;
   16993: out<=0;
   16994: out<=1;
   16995: out<=0;
   16996: out<=1;
   16997: out<=1;
   16998: out<=0;
   16999: out<=0;
   17000: out<=1;
   17001: out<=1;
   17002: out<=1;
   17003: out<=1;
   17004: out<=1;
   17005: out<=0;
   17006: out<=0;
   17007: out<=1;
   17008: out<=1;
   17009: out<=0;
   17010: out<=1;
   17011: out<=0;
   17012: out<=1;
   17013: out<=1;
   17014: out<=0;
   17015: out<=0;
   17016: out<=1;
   17017: out<=1;
   17018: out<=1;
   17019: out<=1;
   17020: out<=1;
   17021: out<=0;
   17022: out<=0;
   17023: out<=1;
   17024: out<=0;
   17025: out<=1;
   17026: out<=0;
   17027: out<=1;
   17028: out<=0;
   17029: out<=0;
   17030: out<=1;
   17031: out<=1;
   17032: out<=0;
   17033: out<=0;
   17034: out<=0;
   17035: out<=0;
   17036: out<=0;
   17037: out<=1;
   17038: out<=1;
   17039: out<=0;
   17040: out<=0;
   17041: out<=1;
   17042: out<=0;
   17043: out<=1;
   17044: out<=0;
   17045: out<=0;
   17046: out<=1;
   17047: out<=1;
   17048: out<=0;
   17049: out<=0;
   17050: out<=0;
   17051: out<=0;
   17052: out<=0;
   17053: out<=1;
   17054: out<=1;
   17055: out<=0;
   17056: out<=1;
   17057: out<=0;
   17058: out<=1;
   17059: out<=0;
   17060: out<=1;
   17061: out<=1;
   17062: out<=0;
   17063: out<=0;
   17064: out<=1;
   17065: out<=1;
   17066: out<=1;
   17067: out<=1;
   17068: out<=1;
   17069: out<=0;
   17070: out<=0;
   17071: out<=1;
   17072: out<=1;
   17073: out<=0;
   17074: out<=1;
   17075: out<=0;
   17076: out<=1;
   17077: out<=1;
   17078: out<=0;
   17079: out<=0;
   17080: out<=1;
   17081: out<=1;
   17082: out<=1;
   17083: out<=1;
   17084: out<=1;
   17085: out<=0;
   17086: out<=0;
   17087: out<=1;
   17088: out<=1;
   17089: out<=0;
   17090: out<=1;
   17091: out<=0;
   17092: out<=1;
   17093: out<=1;
   17094: out<=0;
   17095: out<=0;
   17096: out<=1;
   17097: out<=1;
   17098: out<=1;
   17099: out<=1;
   17100: out<=1;
   17101: out<=0;
   17102: out<=0;
   17103: out<=1;
   17104: out<=0;
   17105: out<=1;
   17106: out<=0;
   17107: out<=1;
   17108: out<=0;
   17109: out<=0;
   17110: out<=1;
   17111: out<=1;
   17112: out<=0;
   17113: out<=0;
   17114: out<=0;
   17115: out<=0;
   17116: out<=0;
   17117: out<=1;
   17118: out<=1;
   17119: out<=0;
   17120: out<=1;
   17121: out<=0;
   17122: out<=1;
   17123: out<=0;
   17124: out<=1;
   17125: out<=1;
   17126: out<=0;
   17127: out<=0;
   17128: out<=1;
   17129: out<=1;
   17130: out<=1;
   17131: out<=1;
   17132: out<=1;
   17133: out<=0;
   17134: out<=0;
   17135: out<=1;
   17136: out<=0;
   17137: out<=1;
   17138: out<=0;
   17139: out<=1;
   17140: out<=0;
   17141: out<=0;
   17142: out<=1;
   17143: out<=1;
   17144: out<=0;
   17145: out<=0;
   17146: out<=0;
   17147: out<=0;
   17148: out<=0;
   17149: out<=1;
   17150: out<=1;
   17151: out<=0;
   17152: out<=0;
   17153: out<=0;
   17154: out<=1;
   17155: out<=1;
   17156: out<=1;
   17157: out<=0;
   17158: out<=1;
   17159: out<=0;
   17160: out<=1;
   17161: out<=0;
   17162: out<=0;
   17163: out<=1;
   17164: out<=0;
   17165: out<=0;
   17166: out<=0;
   17167: out<=0;
   17168: out<=0;
   17169: out<=0;
   17170: out<=1;
   17171: out<=1;
   17172: out<=1;
   17173: out<=0;
   17174: out<=1;
   17175: out<=0;
   17176: out<=1;
   17177: out<=0;
   17178: out<=0;
   17179: out<=1;
   17180: out<=0;
   17181: out<=0;
   17182: out<=0;
   17183: out<=0;
   17184: out<=0;
   17185: out<=0;
   17186: out<=1;
   17187: out<=1;
   17188: out<=1;
   17189: out<=0;
   17190: out<=1;
   17191: out<=0;
   17192: out<=1;
   17193: out<=0;
   17194: out<=0;
   17195: out<=1;
   17196: out<=0;
   17197: out<=0;
   17198: out<=0;
   17199: out<=0;
   17200: out<=0;
   17201: out<=0;
   17202: out<=1;
   17203: out<=1;
   17204: out<=1;
   17205: out<=0;
   17206: out<=1;
   17207: out<=0;
   17208: out<=1;
   17209: out<=0;
   17210: out<=0;
   17211: out<=1;
   17212: out<=0;
   17213: out<=0;
   17214: out<=0;
   17215: out<=0;
   17216: out<=1;
   17217: out<=1;
   17218: out<=0;
   17219: out<=0;
   17220: out<=0;
   17221: out<=1;
   17222: out<=0;
   17223: out<=1;
   17224: out<=0;
   17225: out<=1;
   17226: out<=1;
   17227: out<=0;
   17228: out<=1;
   17229: out<=1;
   17230: out<=1;
   17231: out<=1;
   17232: out<=0;
   17233: out<=0;
   17234: out<=1;
   17235: out<=1;
   17236: out<=1;
   17237: out<=0;
   17238: out<=1;
   17239: out<=0;
   17240: out<=1;
   17241: out<=0;
   17242: out<=0;
   17243: out<=1;
   17244: out<=0;
   17245: out<=0;
   17246: out<=0;
   17247: out<=0;
   17248: out<=0;
   17249: out<=0;
   17250: out<=1;
   17251: out<=1;
   17252: out<=1;
   17253: out<=0;
   17254: out<=1;
   17255: out<=0;
   17256: out<=1;
   17257: out<=0;
   17258: out<=0;
   17259: out<=1;
   17260: out<=0;
   17261: out<=0;
   17262: out<=0;
   17263: out<=0;
   17264: out<=1;
   17265: out<=1;
   17266: out<=0;
   17267: out<=0;
   17268: out<=0;
   17269: out<=1;
   17270: out<=0;
   17271: out<=1;
   17272: out<=0;
   17273: out<=1;
   17274: out<=1;
   17275: out<=0;
   17276: out<=1;
   17277: out<=1;
   17278: out<=1;
   17279: out<=1;
   17280: out<=0;
   17281: out<=0;
   17282: out<=1;
   17283: out<=1;
   17284: out<=1;
   17285: out<=0;
   17286: out<=1;
   17287: out<=0;
   17288: out<=1;
   17289: out<=0;
   17290: out<=0;
   17291: out<=1;
   17292: out<=0;
   17293: out<=0;
   17294: out<=0;
   17295: out<=0;
   17296: out<=1;
   17297: out<=1;
   17298: out<=0;
   17299: out<=0;
   17300: out<=0;
   17301: out<=1;
   17302: out<=0;
   17303: out<=1;
   17304: out<=0;
   17305: out<=1;
   17306: out<=1;
   17307: out<=0;
   17308: out<=1;
   17309: out<=1;
   17310: out<=1;
   17311: out<=1;
   17312: out<=0;
   17313: out<=0;
   17314: out<=1;
   17315: out<=1;
   17316: out<=1;
   17317: out<=0;
   17318: out<=1;
   17319: out<=0;
   17320: out<=1;
   17321: out<=0;
   17322: out<=0;
   17323: out<=1;
   17324: out<=0;
   17325: out<=0;
   17326: out<=0;
   17327: out<=0;
   17328: out<=1;
   17329: out<=1;
   17330: out<=0;
   17331: out<=0;
   17332: out<=0;
   17333: out<=1;
   17334: out<=0;
   17335: out<=1;
   17336: out<=0;
   17337: out<=1;
   17338: out<=1;
   17339: out<=0;
   17340: out<=1;
   17341: out<=1;
   17342: out<=1;
   17343: out<=1;
   17344: out<=1;
   17345: out<=1;
   17346: out<=0;
   17347: out<=0;
   17348: out<=0;
   17349: out<=1;
   17350: out<=0;
   17351: out<=1;
   17352: out<=0;
   17353: out<=1;
   17354: out<=1;
   17355: out<=0;
   17356: out<=1;
   17357: out<=1;
   17358: out<=1;
   17359: out<=1;
   17360: out<=1;
   17361: out<=1;
   17362: out<=0;
   17363: out<=0;
   17364: out<=0;
   17365: out<=1;
   17366: out<=0;
   17367: out<=1;
   17368: out<=0;
   17369: out<=1;
   17370: out<=1;
   17371: out<=0;
   17372: out<=1;
   17373: out<=1;
   17374: out<=1;
   17375: out<=1;
   17376: out<=0;
   17377: out<=0;
   17378: out<=1;
   17379: out<=1;
   17380: out<=1;
   17381: out<=0;
   17382: out<=1;
   17383: out<=0;
   17384: out<=1;
   17385: out<=0;
   17386: out<=0;
   17387: out<=1;
   17388: out<=0;
   17389: out<=0;
   17390: out<=0;
   17391: out<=0;
   17392: out<=0;
   17393: out<=0;
   17394: out<=1;
   17395: out<=1;
   17396: out<=1;
   17397: out<=0;
   17398: out<=1;
   17399: out<=0;
   17400: out<=1;
   17401: out<=0;
   17402: out<=0;
   17403: out<=1;
   17404: out<=0;
   17405: out<=0;
   17406: out<=0;
   17407: out<=0;
   17408: out<=0;
   17409: out<=1;
   17410: out<=1;
   17411: out<=0;
   17412: out<=1;
   17413: out<=1;
   17414: out<=1;
   17415: out<=1;
   17416: out<=0;
   17417: out<=0;
   17418: out<=1;
   17419: out<=1;
   17420: out<=1;
   17421: out<=0;
   17422: out<=1;
   17423: out<=0;
   17424: out<=0;
   17425: out<=1;
   17426: out<=1;
   17427: out<=0;
   17428: out<=1;
   17429: out<=1;
   17430: out<=1;
   17431: out<=1;
   17432: out<=0;
   17433: out<=0;
   17434: out<=1;
   17435: out<=1;
   17436: out<=1;
   17437: out<=0;
   17438: out<=1;
   17439: out<=0;
   17440: out<=1;
   17441: out<=0;
   17442: out<=0;
   17443: out<=1;
   17444: out<=0;
   17445: out<=0;
   17446: out<=0;
   17447: out<=0;
   17448: out<=1;
   17449: out<=1;
   17450: out<=0;
   17451: out<=0;
   17452: out<=0;
   17453: out<=1;
   17454: out<=0;
   17455: out<=1;
   17456: out<=1;
   17457: out<=0;
   17458: out<=0;
   17459: out<=1;
   17460: out<=0;
   17461: out<=0;
   17462: out<=0;
   17463: out<=0;
   17464: out<=1;
   17465: out<=1;
   17466: out<=0;
   17467: out<=0;
   17468: out<=0;
   17469: out<=1;
   17470: out<=0;
   17471: out<=1;
   17472: out<=1;
   17473: out<=0;
   17474: out<=0;
   17475: out<=1;
   17476: out<=0;
   17477: out<=0;
   17478: out<=0;
   17479: out<=0;
   17480: out<=1;
   17481: out<=1;
   17482: out<=0;
   17483: out<=0;
   17484: out<=0;
   17485: out<=1;
   17486: out<=0;
   17487: out<=1;
   17488: out<=0;
   17489: out<=1;
   17490: out<=1;
   17491: out<=0;
   17492: out<=1;
   17493: out<=1;
   17494: out<=1;
   17495: out<=1;
   17496: out<=0;
   17497: out<=0;
   17498: out<=1;
   17499: out<=1;
   17500: out<=1;
   17501: out<=0;
   17502: out<=1;
   17503: out<=0;
   17504: out<=1;
   17505: out<=0;
   17506: out<=0;
   17507: out<=1;
   17508: out<=0;
   17509: out<=0;
   17510: out<=0;
   17511: out<=0;
   17512: out<=1;
   17513: out<=1;
   17514: out<=0;
   17515: out<=0;
   17516: out<=0;
   17517: out<=1;
   17518: out<=0;
   17519: out<=1;
   17520: out<=0;
   17521: out<=1;
   17522: out<=1;
   17523: out<=0;
   17524: out<=1;
   17525: out<=1;
   17526: out<=1;
   17527: out<=1;
   17528: out<=0;
   17529: out<=0;
   17530: out<=1;
   17531: out<=1;
   17532: out<=1;
   17533: out<=0;
   17534: out<=1;
   17535: out<=0;
   17536: out<=0;
   17537: out<=1;
   17538: out<=1;
   17539: out<=0;
   17540: out<=1;
   17541: out<=1;
   17542: out<=1;
   17543: out<=1;
   17544: out<=0;
   17545: out<=0;
   17546: out<=1;
   17547: out<=1;
   17548: out<=1;
   17549: out<=0;
   17550: out<=1;
   17551: out<=0;
   17552: out<=1;
   17553: out<=0;
   17554: out<=0;
   17555: out<=1;
   17556: out<=0;
   17557: out<=0;
   17558: out<=0;
   17559: out<=0;
   17560: out<=1;
   17561: out<=1;
   17562: out<=0;
   17563: out<=0;
   17564: out<=0;
   17565: out<=1;
   17566: out<=0;
   17567: out<=1;
   17568: out<=1;
   17569: out<=0;
   17570: out<=0;
   17571: out<=1;
   17572: out<=0;
   17573: out<=0;
   17574: out<=0;
   17575: out<=0;
   17576: out<=1;
   17577: out<=1;
   17578: out<=0;
   17579: out<=0;
   17580: out<=0;
   17581: out<=1;
   17582: out<=0;
   17583: out<=1;
   17584: out<=0;
   17585: out<=1;
   17586: out<=1;
   17587: out<=0;
   17588: out<=1;
   17589: out<=1;
   17590: out<=1;
   17591: out<=1;
   17592: out<=0;
   17593: out<=0;
   17594: out<=1;
   17595: out<=1;
   17596: out<=1;
   17597: out<=0;
   17598: out<=1;
   17599: out<=0;
   17600: out<=1;
   17601: out<=0;
   17602: out<=0;
   17603: out<=1;
   17604: out<=0;
   17605: out<=0;
   17606: out<=0;
   17607: out<=0;
   17608: out<=1;
   17609: out<=1;
   17610: out<=0;
   17611: out<=0;
   17612: out<=0;
   17613: out<=1;
   17614: out<=0;
   17615: out<=1;
   17616: out<=1;
   17617: out<=0;
   17618: out<=0;
   17619: out<=1;
   17620: out<=0;
   17621: out<=0;
   17622: out<=0;
   17623: out<=0;
   17624: out<=1;
   17625: out<=1;
   17626: out<=0;
   17627: out<=0;
   17628: out<=0;
   17629: out<=1;
   17630: out<=0;
   17631: out<=1;
   17632: out<=1;
   17633: out<=0;
   17634: out<=0;
   17635: out<=1;
   17636: out<=0;
   17637: out<=0;
   17638: out<=0;
   17639: out<=0;
   17640: out<=1;
   17641: out<=1;
   17642: out<=0;
   17643: out<=0;
   17644: out<=0;
   17645: out<=1;
   17646: out<=0;
   17647: out<=1;
   17648: out<=1;
   17649: out<=0;
   17650: out<=0;
   17651: out<=1;
   17652: out<=0;
   17653: out<=0;
   17654: out<=0;
   17655: out<=0;
   17656: out<=1;
   17657: out<=1;
   17658: out<=0;
   17659: out<=0;
   17660: out<=0;
   17661: out<=1;
   17662: out<=0;
   17663: out<=1;
   17664: out<=1;
   17665: out<=1;
   17666: out<=1;
   17667: out<=1;
   17668: out<=1;
   17669: out<=0;
   17670: out<=0;
   17671: out<=1;
   17672: out<=0;
   17673: out<=1;
   17674: out<=0;
   17675: out<=1;
   17676: out<=0;
   17677: out<=0;
   17678: out<=1;
   17679: out<=1;
   17680: out<=0;
   17681: out<=0;
   17682: out<=0;
   17683: out<=0;
   17684: out<=0;
   17685: out<=1;
   17686: out<=1;
   17687: out<=0;
   17688: out<=1;
   17689: out<=0;
   17690: out<=1;
   17691: out<=0;
   17692: out<=1;
   17693: out<=1;
   17694: out<=0;
   17695: out<=0;
   17696: out<=1;
   17697: out<=1;
   17698: out<=1;
   17699: out<=1;
   17700: out<=1;
   17701: out<=0;
   17702: out<=0;
   17703: out<=1;
   17704: out<=0;
   17705: out<=1;
   17706: out<=0;
   17707: out<=1;
   17708: out<=0;
   17709: out<=0;
   17710: out<=1;
   17711: out<=1;
   17712: out<=0;
   17713: out<=0;
   17714: out<=0;
   17715: out<=0;
   17716: out<=0;
   17717: out<=1;
   17718: out<=1;
   17719: out<=0;
   17720: out<=1;
   17721: out<=0;
   17722: out<=1;
   17723: out<=0;
   17724: out<=1;
   17725: out<=1;
   17726: out<=0;
   17727: out<=0;
   17728: out<=0;
   17729: out<=0;
   17730: out<=0;
   17731: out<=0;
   17732: out<=0;
   17733: out<=1;
   17734: out<=1;
   17735: out<=0;
   17736: out<=1;
   17737: out<=0;
   17738: out<=1;
   17739: out<=0;
   17740: out<=1;
   17741: out<=1;
   17742: out<=0;
   17743: out<=0;
   17744: out<=0;
   17745: out<=0;
   17746: out<=0;
   17747: out<=0;
   17748: out<=0;
   17749: out<=1;
   17750: out<=1;
   17751: out<=0;
   17752: out<=1;
   17753: out<=0;
   17754: out<=1;
   17755: out<=0;
   17756: out<=1;
   17757: out<=1;
   17758: out<=0;
   17759: out<=0;
   17760: out<=1;
   17761: out<=1;
   17762: out<=1;
   17763: out<=1;
   17764: out<=1;
   17765: out<=0;
   17766: out<=0;
   17767: out<=1;
   17768: out<=0;
   17769: out<=1;
   17770: out<=0;
   17771: out<=1;
   17772: out<=0;
   17773: out<=0;
   17774: out<=1;
   17775: out<=1;
   17776: out<=1;
   17777: out<=1;
   17778: out<=1;
   17779: out<=1;
   17780: out<=1;
   17781: out<=0;
   17782: out<=0;
   17783: out<=1;
   17784: out<=0;
   17785: out<=1;
   17786: out<=0;
   17787: out<=1;
   17788: out<=0;
   17789: out<=0;
   17790: out<=1;
   17791: out<=1;
   17792: out<=1;
   17793: out<=1;
   17794: out<=1;
   17795: out<=1;
   17796: out<=1;
   17797: out<=0;
   17798: out<=0;
   17799: out<=1;
   17800: out<=0;
   17801: out<=1;
   17802: out<=0;
   17803: out<=1;
   17804: out<=0;
   17805: out<=0;
   17806: out<=1;
   17807: out<=1;
   17808: out<=1;
   17809: out<=1;
   17810: out<=1;
   17811: out<=1;
   17812: out<=1;
   17813: out<=0;
   17814: out<=0;
   17815: out<=1;
   17816: out<=0;
   17817: out<=1;
   17818: out<=0;
   17819: out<=1;
   17820: out<=0;
   17821: out<=0;
   17822: out<=1;
   17823: out<=1;
   17824: out<=1;
   17825: out<=1;
   17826: out<=1;
   17827: out<=1;
   17828: out<=1;
   17829: out<=0;
   17830: out<=0;
   17831: out<=1;
   17832: out<=0;
   17833: out<=1;
   17834: out<=0;
   17835: out<=1;
   17836: out<=0;
   17837: out<=0;
   17838: out<=1;
   17839: out<=1;
   17840: out<=1;
   17841: out<=1;
   17842: out<=1;
   17843: out<=1;
   17844: out<=1;
   17845: out<=0;
   17846: out<=0;
   17847: out<=1;
   17848: out<=0;
   17849: out<=1;
   17850: out<=0;
   17851: out<=1;
   17852: out<=0;
   17853: out<=0;
   17854: out<=1;
   17855: out<=1;
   17856: out<=0;
   17857: out<=0;
   17858: out<=0;
   17859: out<=0;
   17860: out<=0;
   17861: out<=1;
   17862: out<=1;
   17863: out<=0;
   17864: out<=1;
   17865: out<=0;
   17866: out<=1;
   17867: out<=0;
   17868: out<=1;
   17869: out<=1;
   17870: out<=0;
   17871: out<=0;
   17872: out<=1;
   17873: out<=1;
   17874: out<=1;
   17875: out<=1;
   17876: out<=1;
   17877: out<=0;
   17878: out<=0;
   17879: out<=1;
   17880: out<=0;
   17881: out<=1;
   17882: out<=0;
   17883: out<=1;
   17884: out<=0;
   17885: out<=0;
   17886: out<=1;
   17887: out<=1;
   17888: out<=1;
   17889: out<=1;
   17890: out<=1;
   17891: out<=1;
   17892: out<=1;
   17893: out<=0;
   17894: out<=0;
   17895: out<=1;
   17896: out<=0;
   17897: out<=1;
   17898: out<=0;
   17899: out<=1;
   17900: out<=0;
   17901: out<=0;
   17902: out<=1;
   17903: out<=1;
   17904: out<=0;
   17905: out<=0;
   17906: out<=0;
   17907: out<=0;
   17908: out<=0;
   17909: out<=1;
   17910: out<=1;
   17911: out<=0;
   17912: out<=1;
   17913: out<=0;
   17914: out<=1;
   17915: out<=0;
   17916: out<=1;
   17917: out<=1;
   17918: out<=0;
   17919: out<=0;
   17920: out<=1;
   17921: out<=1;
   17922: out<=0;
   17923: out<=0;
   17924: out<=1;
   17925: out<=0;
   17926: out<=1;
   17927: out<=0;
   17928: out<=1;
   17929: out<=0;
   17930: out<=0;
   17931: out<=1;
   17932: out<=1;
   17933: out<=1;
   17934: out<=1;
   17935: out<=1;
   17936: out<=0;
   17937: out<=0;
   17938: out<=1;
   17939: out<=1;
   17940: out<=0;
   17941: out<=1;
   17942: out<=0;
   17943: out<=1;
   17944: out<=0;
   17945: out<=1;
   17946: out<=1;
   17947: out<=0;
   17948: out<=0;
   17949: out<=0;
   17950: out<=0;
   17951: out<=0;
   17952: out<=0;
   17953: out<=0;
   17954: out<=1;
   17955: out<=1;
   17956: out<=0;
   17957: out<=1;
   17958: out<=0;
   17959: out<=1;
   17960: out<=0;
   17961: out<=1;
   17962: out<=1;
   17963: out<=0;
   17964: out<=0;
   17965: out<=0;
   17966: out<=0;
   17967: out<=0;
   17968: out<=1;
   17969: out<=1;
   17970: out<=0;
   17971: out<=0;
   17972: out<=1;
   17973: out<=0;
   17974: out<=1;
   17975: out<=0;
   17976: out<=1;
   17977: out<=0;
   17978: out<=0;
   17979: out<=1;
   17980: out<=1;
   17981: out<=1;
   17982: out<=1;
   17983: out<=1;
   17984: out<=0;
   17985: out<=0;
   17986: out<=1;
   17987: out<=1;
   17988: out<=0;
   17989: out<=1;
   17990: out<=0;
   17991: out<=1;
   17992: out<=0;
   17993: out<=1;
   17994: out<=1;
   17995: out<=0;
   17996: out<=0;
   17997: out<=0;
   17998: out<=0;
   17999: out<=0;
   18000: out<=0;
   18001: out<=0;
   18002: out<=1;
   18003: out<=1;
   18004: out<=0;
   18005: out<=1;
   18006: out<=0;
   18007: out<=1;
   18008: out<=0;
   18009: out<=1;
   18010: out<=1;
   18011: out<=0;
   18012: out<=0;
   18013: out<=0;
   18014: out<=0;
   18015: out<=0;
   18016: out<=0;
   18017: out<=0;
   18018: out<=1;
   18019: out<=1;
   18020: out<=0;
   18021: out<=1;
   18022: out<=0;
   18023: out<=1;
   18024: out<=0;
   18025: out<=1;
   18026: out<=1;
   18027: out<=0;
   18028: out<=0;
   18029: out<=0;
   18030: out<=0;
   18031: out<=0;
   18032: out<=0;
   18033: out<=0;
   18034: out<=1;
   18035: out<=1;
   18036: out<=0;
   18037: out<=1;
   18038: out<=0;
   18039: out<=1;
   18040: out<=0;
   18041: out<=1;
   18042: out<=1;
   18043: out<=0;
   18044: out<=0;
   18045: out<=0;
   18046: out<=0;
   18047: out<=0;
   18048: out<=1;
   18049: out<=1;
   18050: out<=0;
   18051: out<=0;
   18052: out<=1;
   18053: out<=0;
   18054: out<=1;
   18055: out<=0;
   18056: out<=1;
   18057: out<=0;
   18058: out<=0;
   18059: out<=1;
   18060: out<=1;
   18061: out<=1;
   18062: out<=1;
   18063: out<=1;
   18064: out<=1;
   18065: out<=1;
   18066: out<=0;
   18067: out<=0;
   18068: out<=1;
   18069: out<=0;
   18070: out<=1;
   18071: out<=0;
   18072: out<=1;
   18073: out<=0;
   18074: out<=0;
   18075: out<=1;
   18076: out<=1;
   18077: out<=1;
   18078: out<=1;
   18079: out<=1;
   18080: out<=0;
   18081: out<=0;
   18082: out<=1;
   18083: out<=1;
   18084: out<=0;
   18085: out<=1;
   18086: out<=0;
   18087: out<=1;
   18088: out<=0;
   18089: out<=1;
   18090: out<=1;
   18091: out<=0;
   18092: out<=0;
   18093: out<=0;
   18094: out<=0;
   18095: out<=0;
   18096: out<=0;
   18097: out<=0;
   18098: out<=1;
   18099: out<=1;
   18100: out<=0;
   18101: out<=1;
   18102: out<=0;
   18103: out<=1;
   18104: out<=0;
   18105: out<=1;
   18106: out<=1;
   18107: out<=0;
   18108: out<=0;
   18109: out<=0;
   18110: out<=0;
   18111: out<=0;
   18112: out<=0;
   18113: out<=0;
   18114: out<=1;
   18115: out<=1;
   18116: out<=0;
   18117: out<=1;
   18118: out<=0;
   18119: out<=1;
   18120: out<=0;
   18121: out<=1;
   18122: out<=1;
   18123: out<=0;
   18124: out<=0;
   18125: out<=0;
   18126: out<=0;
   18127: out<=0;
   18128: out<=1;
   18129: out<=1;
   18130: out<=0;
   18131: out<=0;
   18132: out<=1;
   18133: out<=0;
   18134: out<=1;
   18135: out<=0;
   18136: out<=1;
   18137: out<=0;
   18138: out<=0;
   18139: out<=1;
   18140: out<=1;
   18141: out<=1;
   18142: out<=1;
   18143: out<=1;
   18144: out<=0;
   18145: out<=0;
   18146: out<=1;
   18147: out<=1;
   18148: out<=0;
   18149: out<=1;
   18150: out<=0;
   18151: out<=1;
   18152: out<=0;
   18153: out<=1;
   18154: out<=1;
   18155: out<=0;
   18156: out<=0;
   18157: out<=0;
   18158: out<=0;
   18159: out<=0;
   18160: out<=1;
   18161: out<=1;
   18162: out<=0;
   18163: out<=0;
   18164: out<=1;
   18165: out<=0;
   18166: out<=1;
   18167: out<=0;
   18168: out<=1;
   18169: out<=0;
   18170: out<=0;
   18171: out<=1;
   18172: out<=1;
   18173: out<=1;
   18174: out<=1;
   18175: out<=1;
   18176: out<=0;
   18177: out<=1;
   18178: out<=0;
   18179: out<=1;
   18180: out<=1;
   18181: out<=1;
   18182: out<=0;
   18183: out<=0;
   18184: out<=1;
   18185: out<=1;
   18186: out<=1;
   18187: out<=1;
   18188: out<=0;
   18189: out<=1;
   18190: out<=1;
   18191: out<=0;
   18192: out<=0;
   18193: out<=1;
   18194: out<=0;
   18195: out<=1;
   18196: out<=1;
   18197: out<=1;
   18198: out<=0;
   18199: out<=0;
   18200: out<=1;
   18201: out<=1;
   18202: out<=1;
   18203: out<=1;
   18204: out<=0;
   18205: out<=1;
   18206: out<=1;
   18207: out<=0;
   18208: out<=0;
   18209: out<=1;
   18210: out<=0;
   18211: out<=1;
   18212: out<=1;
   18213: out<=1;
   18214: out<=0;
   18215: out<=0;
   18216: out<=1;
   18217: out<=1;
   18218: out<=1;
   18219: out<=1;
   18220: out<=0;
   18221: out<=1;
   18222: out<=1;
   18223: out<=0;
   18224: out<=0;
   18225: out<=1;
   18226: out<=0;
   18227: out<=1;
   18228: out<=1;
   18229: out<=1;
   18230: out<=0;
   18231: out<=0;
   18232: out<=1;
   18233: out<=1;
   18234: out<=1;
   18235: out<=1;
   18236: out<=0;
   18237: out<=1;
   18238: out<=1;
   18239: out<=0;
   18240: out<=1;
   18241: out<=0;
   18242: out<=1;
   18243: out<=0;
   18244: out<=0;
   18245: out<=0;
   18246: out<=1;
   18247: out<=1;
   18248: out<=0;
   18249: out<=0;
   18250: out<=0;
   18251: out<=0;
   18252: out<=1;
   18253: out<=0;
   18254: out<=0;
   18255: out<=1;
   18256: out<=0;
   18257: out<=1;
   18258: out<=0;
   18259: out<=1;
   18260: out<=1;
   18261: out<=1;
   18262: out<=0;
   18263: out<=0;
   18264: out<=1;
   18265: out<=1;
   18266: out<=1;
   18267: out<=1;
   18268: out<=0;
   18269: out<=1;
   18270: out<=1;
   18271: out<=0;
   18272: out<=0;
   18273: out<=1;
   18274: out<=0;
   18275: out<=1;
   18276: out<=1;
   18277: out<=1;
   18278: out<=0;
   18279: out<=0;
   18280: out<=1;
   18281: out<=1;
   18282: out<=1;
   18283: out<=1;
   18284: out<=0;
   18285: out<=1;
   18286: out<=1;
   18287: out<=0;
   18288: out<=1;
   18289: out<=0;
   18290: out<=1;
   18291: out<=0;
   18292: out<=0;
   18293: out<=0;
   18294: out<=1;
   18295: out<=1;
   18296: out<=0;
   18297: out<=0;
   18298: out<=0;
   18299: out<=0;
   18300: out<=1;
   18301: out<=0;
   18302: out<=0;
   18303: out<=1;
   18304: out<=0;
   18305: out<=1;
   18306: out<=0;
   18307: out<=1;
   18308: out<=1;
   18309: out<=1;
   18310: out<=0;
   18311: out<=0;
   18312: out<=1;
   18313: out<=1;
   18314: out<=1;
   18315: out<=1;
   18316: out<=0;
   18317: out<=1;
   18318: out<=1;
   18319: out<=0;
   18320: out<=1;
   18321: out<=0;
   18322: out<=1;
   18323: out<=0;
   18324: out<=0;
   18325: out<=0;
   18326: out<=1;
   18327: out<=1;
   18328: out<=0;
   18329: out<=0;
   18330: out<=0;
   18331: out<=0;
   18332: out<=1;
   18333: out<=0;
   18334: out<=0;
   18335: out<=1;
   18336: out<=0;
   18337: out<=1;
   18338: out<=0;
   18339: out<=1;
   18340: out<=1;
   18341: out<=1;
   18342: out<=0;
   18343: out<=0;
   18344: out<=1;
   18345: out<=1;
   18346: out<=1;
   18347: out<=1;
   18348: out<=0;
   18349: out<=1;
   18350: out<=1;
   18351: out<=0;
   18352: out<=1;
   18353: out<=0;
   18354: out<=1;
   18355: out<=0;
   18356: out<=0;
   18357: out<=0;
   18358: out<=1;
   18359: out<=1;
   18360: out<=0;
   18361: out<=0;
   18362: out<=0;
   18363: out<=0;
   18364: out<=1;
   18365: out<=0;
   18366: out<=0;
   18367: out<=1;
   18368: out<=1;
   18369: out<=0;
   18370: out<=1;
   18371: out<=0;
   18372: out<=0;
   18373: out<=0;
   18374: out<=1;
   18375: out<=1;
   18376: out<=0;
   18377: out<=0;
   18378: out<=0;
   18379: out<=0;
   18380: out<=1;
   18381: out<=0;
   18382: out<=0;
   18383: out<=1;
   18384: out<=1;
   18385: out<=0;
   18386: out<=1;
   18387: out<=0;
   18388: out<=0;
   18389: out<=0;
   18390: out<=1;
   18391: out<=1;
   18392: out<=0;
   18393: out<=0;
   18394: out<=0;
   18395: out<=0;
   18396: out<=1;
   18397: out<=0;
   18398: out<=0;
   18399: out<=1;
   18400: out<=0;
   18401: out<=1;
   18402: out<=0;
   18403: out<=1;
   18404: out<=1;
   18405: out<=1;
   18406: out<=0;
   18407: out<=0;
   18408: out<=1;
   18409: out<=1;
   18410: out<=1;
   18411: out<=1;
   18412: out<=0;
   18413: out<=1;
   18414: out<=1;
   18415: out<=0;
   18416: out<=0;
   18417: out<=1;
   18418: out<=0;
   18419: out<=1;
   18420: out<=1;
   18421: out<=1;
   18422: out<=0;
   18423: out<=0;
   18424: out<=1;
   18425: out<=1;
   18426: out<=1;
   18427: out<=1;
   18428: out<=0;
   18429: out<=1;
   18430: out<=1;
   18431: out<=0;
   18432: out<=0;
   18433: out<=1;
   18434: out<=0;
   18435: out<=1;
   18436: out<=1;
   18437: out<=1;
   18438: out<=0;
   18439: out<=0;
   18440: out<=0;
   18441: out<=0;
   18442: out<=0;
   18443: out<=0;
   18444: out<=1;
   18445: out<=0;
   18446: out<=0;
   18447: out<=1;
   18448: out<=0;
   18449: out<=1;
   18450: out<=0;
   18451: out<=1;
   18452: out<=1;
   18453: out<=1;
   18454: out<=0;
   18455: out<=0;
   18456: out<=0;
   18457: out<=0;
   18458: out<=0;
   18459: out<=0;
   18460: out<=1;
   18461: out<=0;
   18462: out<=0;
   18463: out<=1;
   18464: out<=1;
   18465: out<=0;
   18466: out<=1;
   18467: out<=0;
   18468: out<=0;
   18469: out<=0;
   18470: out<=1;
   18471: out<=1;
   18472: out<=1;
   18473: out<=1;
   18474: out<=1;
   18475: out<=1;
   18476: out<=0;
   18477: out<=1;
   18478: out<=1;
   18479: out<=0;
   18480: out<=1;
   18481: out<=0;
   18482: out<=1;
   18483: out<=0;
   18484: out<=0;
   18485: out<=0;
   18486: out<=1;
   18487: out<=1;
   18488: out<=1;
   18489: out<=1;
   18490: out<=1;
   18491: out<=1;
   18492: out<=0;
   18493: out<=1;
   18494: out<=1;
   18495: out<=0;
   18496: out<=1;
   18497: out<=0;
   18498: out<=1;
   18499: out<=0;
   18500: out<=0;
   18501: out<=0;
   18502: out<=1;
   18503: out<=1;
   18504: out<=1;
   18505: out<=1;
   18506: out<=1;
   18507: out<=1;
   18508: out<=0;
   18509: out<=1;
   18510: out<=1;
   18511: out<=0;
   18512: out<=0;
   18513: out<=1;
   18514: out<=0;
   18515: out<=1;
   18516: out<=1;
   18517: out<=1;
   18518: out<=0;
   18519: out<=0;
   18520: out<=0;
   18521: out<=0;
   18522: out<=0;
   18523: out<=0;
   18524: out<=1;
   18525: out<=0;
   18526: out<=0;
   18527: out<=1;
   18528: out<=1;
   18529: out<=0;
   18530: out<=1;
   18531: out<=0;
   18532: out<=0;
   18533: out<=0;
   18534: out<=1;
   18535: out<=1;
   18536: out<=1;
   18537: out<=1;
   18538: out<=1;
   18539: out<=1;
   18540: out<=0;
   18541: out<=1;
   18542: out<=1;
   18543: out<=0;
   18544: out<=0;
   18545: out<=1;
   18546: out<=0;
   18547: out<=1;
   18548: out<=1;
   18549: out<=1;
   18550: out<=0;
   18551: out<=0;
   18552: out<=0;
   18553: out<=0;
   18554: out<=0;
   18555: out<=0;
   18556: out<=1;
   18557: out<=0;
   18558: out<=0;
   18559: out<=1;
   18560: out<=0;
   18561: out<=1;
   18562: out<=0;
   18563: out<=1;
   18564: out<=1;
   18565: out<=1;
   18566: out<=0;
   18567: out<=0;
   18568: out<=0;
   18569: out<=0;
   18570: out<=0;
   18571: out<=0;
   18572: out<=1;
   18573: out<=0;
   18574: out<=0;
   18575: out<=1;
   18576: out<=1;
   18577: out<=0;
   18578: out<=1;
   18579: out<=0;
   18580: out<=0;
   18581: out<=0;
   18582: out<=1;
   18583: out<=1;
   18584: out<=1;
   18585: out<=1;
   18586: out<=1;
   18587: out<=1;
   18588: out<=0;
   18589: out<=1;
   18590: out<=1;
   18591: out<=0;
   18592: out<=1;
   18593: out<=0;
   18594: out<=1;
   18595: out<=0;
   18596: out<=0;
   18597: out<=0;
   18598: out<=1;
   18599: out<=1;
   18600: out<=1;
   18601: out<=1;
   18602: out<=1;
   18603: out<=1;
   18604: out<=0;
   18605: out<=1;
   18606: out<=1;
   18607: out<=0;
   18608: out<=0;
   18609: out<=1;
   18610: out<=0;
   18611: out<=1;
   18612: out<=1;
   18613: out<=1;
   18614: out<=0;
   18615: out<=0;
   18616: out<=0;
   18617: out<=0;
   18618: out<=0;
   18619: out<=0;
   18620: out<=1;
   18621: out<=0;
   18622: out<=0;
   18623: out<=1;
   18624: out<=1;
   18625: out<=0;
   18626: out<=1;
   18627: out<=0;
   18628: out<=0;
   18629: out<=0;
   18630: out<=1;
   18631: out<=1;
   18632: out<=1;
   18633: out<=1;
   18634: out<=1;
   18635: out<=1;
   18636: out<=0;
   18637: out<=1;
   18638: out<=1;
   18639: out<=0;
   18640: out<=1;
   18641: out<=0;
   18642: out<=1;
   18643: out<=0;
   18644: out<=0;
   18645: out<=0;
   18646: out<=1;
   18647: out<=1;
   18648: out<=1;
   18649: out<=1;
   18650: out<=1;
   18651: out<=1;
   18652: out<=0;
   18653: out<=1;
   18654: out<=1;
   18655: out<=0;
   18656: out<=1;
   18657: out<=0;
   18658: out<=1;
   18659: out<=0;
   18660: out<=0;
   18661: out<=0;
   18662: out<=1;
   18663: out<=1;
   18664: out<=1;
   18665: out<=1;
   18666: out<=1;
   18667: out<=1;
   18668: out<=0;
   18669: out<=1;
   18670: out<=1;
   18671: out<=0;
   18672: out<=1;
   18673: out<=0;
   18674: out<=1;
   18675: out<=0;
   18676: out<=0;
   18677: out<=0;
   18678: out<=1;
   18679: out<=1;
   18680: out<=1;
   18681: out<=1;
   18682: out<=1;
   18683: out<=1;
   18684: out<=0;
   18685: out<=1;
   18686: out<=1;
   18687: out<=0;
   18688: out<=1;
   18689: out<=1;
   18690: out<=0;
   18691: out<=0;
   18692: out<=1;
   18693: out<=0;
   18694: out<=1;
   18695: out<=0;
   18696: out<=0;
   18697: out<=1;
   18698: out<=1;
   18699: out<=0;
   18700: out<=0;
   18701: out<=0;
   18702: out<=0;
   18703: out<=0;
   18704: out<=0;
   18705: out<=0;
   18706: out<=1;
   18707: out<=1;
   18708: out<=0;
   18709: out<=1;
   18710: out<=0;
   18711: out<=1;
   18712: out<=1;
   18713: out<=0;
   18714: out<=0;
   18715: out<=1;
   18716: out<=1;
   18717: out<=1;
   18718: out<=1;
   18719: out<=1;
   18720: out<=1;
   18721: out<=1;
   18722: out<=0;
   18723: out<=0;
   18724: out<=1;
   18725: out<=0;
   18726: out<=1;
   18727: out<=0;
   18728: out<=0;
   18729: out<=1;
   18730: out<=1;
   18731: out<=0;
   18732: out<=0;
   18733: out<=0;
   18734: out<=0;
   18735: out<=0;
   18736: out<=0;
   18737: out<=0;
   18738: out<=1;
   18739: out<=1;
   18740: out<=0;
   18741: out<=1;
   18742: out<=0;
   18743: out<=1;
   18744: out<=1;
   18745: out<=0;
   18746: out<=0;
   18747: out<=1;
   18748: out<=1;
   18749: out<=1;
   18750: out<=1;
   18751: out<=1;
   18752: out<=0;
   18753: out<=0;
   18754: out<=1;
   18755: out<=1;
   18756: out<=0;
   18757: out<=1;
   18758: out<=0;
   18759: out<=1;
   18760: out<=1;
   18761: out<=0;
   18762: out<=0;
   18763: out<=1;
   18764: out<=1;
   18765: out<=1;
   18766: out<=1;
   18767: out<=1;
   18768: out<=0;
   18769: out<=0;
   18770: out<=1;
   18771: out<=1;
   18772: out<=0;
   18773: out<=1;
   18774: out<=0;
   18775: out<=1;
   18776: out<=1;
   18777: out<=0;
   18778: out<=0;
   18779: out<=1;
   18780: out<=1;
   18781: out<=1;
   18782: out<=1;
   18783: out<=1;
   18784: out<=1;
   18785: out<=1;
   18786: out<=0;
   18787: out<=0;
   18788: out<=1;
   18789: out<=0;
   18790: out<=1;
   18791: out<=0;
   18792: out<=0;
   18793: out<=1;
   18794: out<=1;
   18795: out<=0;
   18796: out<=0;
   18797: out<=0;
   18798: out<=0;
   18799: out<=0;
   18800: out<=1;
   18801: out<=1;
   18802: out<=0;
   18803: out<=0;
   18804: out<=1;
   18805: out<=0;
   18806: out<=1;
   18807: out<=0;
   18808: out<=0;
   18809: out<=1;
   18810: out<=1;
   18811: out<=0;
   18812: out<=0;
   18813: out<=0;
   18814: out<=0;
   18815: out<=0;
   18816: out<=1;
   18817: out<=1;
   18818: out<=0;
   18819: out<=0;
   18820: out<=1;
   18821: out<=0;
   18822: out<=1;
   18823: out<=0;
   18824: out<=0;
   18825: out<=1;
   18826: out<=1;
   18827: out<=0;
   18828: out<=0;
   18829: out<=0;
   18830: out<=0;
   18831: out<=0;
   18832: out<=1;
   18833: out<=1;
   18834: out<=0;
   18835: out<=0;
   18836: out<=1;
   18837: out<=0;
   18838: out<=1;
   18839: out<=0;
   18840: out<=0;
   18841: out<=1;
   18842: out<=1;
   18843: out<=0;
   18844: out<=0;
   18845: out<=0;
   18846: out<=0;
   18847: out<=0;
   18848: out<=1;
   18849: out<=1;
   18850: out<=0;
   18851: out<=0;
   18852: out<=1;
   18853: out<=0;
   18854: out<=1;
   18855: out<=0;
   18856: out<=0;
   18857: out<=1;
   18858: out<=1;
   18859: out<=0;
   18860: out<=0;
   18861: out<=0;
   18862: out<=0;
   18863: out<=0;
   18864: out<=1;
   18865: out<=1;
   18866: out<=0;
   18867: out<=0;
   18868: out<=1;
   18869: out<=0;
   18870: out<=1;
   18871: out<=0;
   18872: out<=0;
   18873: out<=1;
   18874: out<=1;
   18875: out<=0;
   18876: out<=0;
   18877: out<=0;
   18878: out<=0;
   18879: out<=0;
   18880: out<=0;
   18881: out<=0;
   18882: out<=1;
   18883: out<=1;
   18884: out<=0;
   18885: out<=1;
   18886: out<=0;
   18887: out<=1;
   18888: out<=1;
   18889: out<=0;
   18890: out<=0;
   18891: out<=1;
   18892: out<=1;
   18893: out<=1;
   18894: out<=1;
   18895: out<=1;
   18896: out<=1;
   18897: out<=1;
   18898: out<=0;
   18899: out<=0;
   18900: out<=1;
   18901: out<=0;
   18902: out<=1;
   18903: out<=0;
   18904: out<=0;
   18905: out<=1;
   18906: out<=1;
   18907: out<=0;
   18908: out<=0;
   18909: out<=0;
   18910: out<=0;
   18911: out<=0;
   18912: out<=1;
   18913: out<=1;
   18914: out<=0;
   18915: out<=0;
   18916: out<=1;
   18917: out<=0;
   18918: out<=1;
   18919: out<=0;
   18920: out<=0;
   18921: out<=1;
   18922: out<=1;
   18923: out<=0;
   18924: out<=0;
   18925: out<=0;
   18926: out<=0;
   18927: out<=0;
   18928: out<=0;
   18929: out<=0;
   18930: out<=1;
   18931: out<=1;
   18932: out<=0;
   18933: out<=1;
   18934: out<=0;
   18935: out<=1;
   18936: out<=1;
   18937: out<=0;
   18938: out<=0;
   18939: out<=1;
   18940: out<=1;
   18941: out<=1;
   18942: out<=1;
   18943: out<=1;
   18944: out<=0;
   18945: out<=0;
   18946: out<=0;
   18947: out<=0;
   18948: out<=0;
   18949: out<=1;
   18950: out<=1;
   18951: out<=0;
   18952: out<=0;
   18953: out<=1;
   18954: out<=0;
   18955: out<=1;
   18956: out<=0;
   18957: out<=0;
   18958: out<=1;
   18959: out<=1;
   18960: out<=1;
   18961: out<=1;
   18962: out<=1;
   18963: out<=1;
   18964: out<=1;
   18965: out<=0;
   18966: out<=0;
   18967: out<=1;
   18968: out<=1;
   18969: out<=0;
   18970: out<=1;
   18971: out<=0;
   18972: out<=1;
   18973: out<=1;
   18974: out<=0;
   18975: out<=0;
   18976: out<=1;
   18977: out<=1;
   18978: out<=1;
   18979: out<=1;
   18980: out<=1;
   18981: out<=0;
   18982: out<=0;
   18983: out<=1;
   18984: out<=1;
   18985: out<=0;
   18986: out<=1;
   18987: out<=0;
   18988: out<=1;
   18989: out<=1;
   18990: out<=0;
   18991: out<=0;
   18992: out<=0;
   18993: out<=0;
   18994: out<=0;
   18995: out<=0;
   18996: out<=0;
   18997: out<=1;
   18998: out<=1;
   18999: out<=0;
   19000: out<=0;
   19001: out<=1;
   19002: out<=0;
   19003: out<=1;
   19004: out<=0;
   19005: out<=0;
   19006: out<=1;
   19007: out<=1;
   19008: out<=1;
   19009: out<=1;
   19010: out<=1;
   19011: out<=1;
   19012: out<=1;
   19013: out<=0;
   19014: out<=0;
   19015: out<=1;
   19016: out<=1;
   19017: out<=0;
   19018: out<=1;
   19019: out<=0;
   19020: out<=1;
   19021: out<=1;
   19022: out<=0;
   19023: out<=0;
   19024: out<=1;
   19025: out<=1;
   19026: out<=1;
   19027: out<=1;
   19028: out<=1;
   19029: out<=0;
   19030: out<=0;
   19031: out<=1;
   19032: out<=1;
   19033: out<=0;
   19034: out<=1;
   19035: out<=0;
   19036: out<=1;
   19037: out<=1;
   19038: out<=0;
   19039: out<=0;
   19040: out<=1;
   19041: out<=1;
   19042: out<=1;
   19043: out<=1;
   19044: out<=1;
   19045: out<=0;
   19046: out<=0;
   19047: out<=1;
   19048: out<=1;
   19049: out<=0;
   19050: out<=1;
   19051: out<=0;
   19052: out<=1;
   19053: out<=1;
   19054: out<=0;
   19055: out<=0;
   19056: out<=1;
   19057: out<=1;
   19058: out<=1;
   19059: out<=1;
   19060: out<=1;
   19061: out<=0;
   19062: out<=0;
   19063: out<=1;
   19064: out<=1;
   19065: out<=0;
   19066: out<=1;
   19067: out<=0;
   19068: out<=1;
   19069: out<=1;
   19070: out<=0;
   19071: out<=0;
   19072: out<=0;
   19073: out<=0;
   19074: out<=0;
   19075: out<=0;
   19076: out<=0;
   19077: out<=1;
   19078: out<=1;
   19079: out<=0;
   19080: out<=0;
   19081: out<=1;
   19082: out<=0;
   19083: out<=1;
   19084: out<=0;
   19085: out<=0;
   19086: out<=1;
   19087: out<=1;
   19088: out<=0;
   19089: out<=0;
   19090: out<=0;
   19091: out<=0;
   19092: out<=0;
   19093: out<=1;
   19094: out<=1;
   19095: out<=0;
   19096: out<=0;
   19097: out<=1;
   19098: out<=0;
   19099: out<=1;
   19100: out<=0;
   19101: out<=0;
   19102: out<=1;
   19103: out<=1;
   19104: out<=1;
   19105: out<=1;
   19106: out<=1;
   19107: out<=1;
   19108: out<=1;
   19109: out<=0;
   19110: out<=0;
   19111: out<=1;
   19112: out<=1;
   19113: out<=0;
   19114: out<=1;
   19115: out<=0;
   19116: out<=1;
   19117: out<=1;
   19118: out<=0;
   19119: out<=0;
   19120: out<=1;
   19121: out<=1;
   19122: out<=1;
   19123: out<=1;
   19124: out<=1;
   19125: out<=0;
   19126: out<=0;
   19127: out<=1;
   19128: out<=1;
   19129: out<=0;
   19130: out<=1;
   19131: out<=0;
   19132: out<=1;
   19133: out<=1;
   19134: out<=0;
   19135: out<=0;
   19136: out<=1;
   19137: out<=1;
   19138: out<=1;
   19139: out<=1;
   19140: out<=1;
   19141: out<=0;
   19142: out<=0;
   19143: out<=1;
   19144: out<=1;
   19145: out<=0;
   19146: out<=1;
   19147: out<=0;
   19148: out<=1;
   19149: out<=1;
   19150: out<=0;
   19151: out<=0;
   19152: out<=0;
   19153: out<=0;
   19154: out<=0;
   19155: out<=0;
   19156: out<=0;
   19157: out<=1;
   19158: out<=1;
   19159: out<=0;
   19160: out<=0;
   19161: out<=1;
   19162: out<=0;
   19163: out<=1;
   19164: out<=0;
   19165: out<=0;
   19166: out<=1;
   19167: out<=1;
   19168: out<=1;
   19169: out<=1;
   19170: out<=1;
   19171: out<=1;
   19172: out<=1;
   19173: out<=0;
   19174: out<=0;
   19175: out<=1;
   19176: out<=1;
   19177: out<=0;
   19178: out<=1;
   19179: out<=0;
   19180: out<=1;
   19181: out<=1;
   19182: out<=0;
   19183: out<=0;
   19184: out<=0;
   19185: out<=0;
   19186: out<=0;
   19187: out<=0;
   19188: out<=0;
   19189: out<=1;
   19190: out<=1;
   19191: out<=0;
   19192: out<=0;
   19193: out<=1;
   19194: out<=0;
   19195: out<=1;
   19196: out<=0;
   19197: out<=0;
   19198: out<=1;
   19199: out<=1;
   19200: out<=1;
   19201: out<=0;
   19202: out<=0;
   19203: out<=1;
   19204: out<=0;
   19205: out<=0;
   19206: out<=0;
   19207: out<=0;
   19208: out<=0;
   19209: out<=0;
   19210: out<=1;
   19211: out<=1;
   19212: out<=1;
   19213: out<=0;
   19214: out<=1;
   19215: out<=0;
   19216: out<=1;
   19217: out<=0;
   19218: out<=0;
   19219: out<=1;
   19220: out<=0;
   19221: out<=0;
   19222: out<=0;
   19223: out<=0;
   19224: out<=0;
   19225: out<=0;
   19226: out<=1;
   19227: out<=1;
   19228: out<=1;
   19229: out<=0;
   19230: out<=1;
   19231: out<=0;
   19232: out<=1;
   19233: out<=0;
   19234: out<=0;
   19235: out<=1;
   19236: out<=0;
   19237: out<=0;
   19238: out<=0;
   19239: out<=0;
   19240: out<=0;
   19241: out<=0;
   19242: out<=1;
   19243: out<=1;
   19244: out<=1;
   19245: out<=0;
   19246: out<=1;
   19247: out<=0;
   19248: out<=1;
   19249: out<=0;
   19250: out<=0;
   19251: out<=1;
   19252: out<=0;
   19253: out<=0;
   19254: out<=0;
   19255: out<=0;
   19256: out<=0;
   19257: out<=0;
   19258: out<=1;
   19259: out<=1;
   19260: out<=1;
   19261: out<=0;
   19262: out<=1;
   19263: out<=0;
   19264: out<=0;
   19265: out<=1;
   19266: out<=1;
   19267: out<=0;
   19268: out<=1;
   19269: out<=1;
   19270: out<=1;
   19271: out<=1;
   19272: out<=1;
   19273: out<=1;
   19274: out<=0;
   19275: out<=0;
   19276: out<=0;
   19277: out<=1;
   19278: out<=0;
   19279: out<=1;
   19280: out<=1;
   19281: out<=0;
   19282: out<=0;
   19283: out<=1;
   19284: out<=0;
   19285: out<=0;
   19286: out<=0;
   19287: out<=0;
   19288: out<=0;
   19289: out<=0;
   19290: out<=1;
   19291: out<=1;
   19292: out<=1;
   19293: out<=0;
   19294: out<=1;
   19295: out<=0;
   19296: out<=1;
   19297: out<=0;
   19298: out<=0;
   19299: out<=1;
   19300: out<=0;
   19301: out<=0;
   19302: out<=0;
   19303: out<=0;
   19304: out<=0;
   19305: out<=0;
   19306: out<=1;
   19307: out<=1;
   19308: out<=1;
   19309: out<=0;
   19310: out<=1;
   19311: out<=0;
   19312: out<=0;
   19313: out<=1;
   19314: out<=1;
   19315: out<=0;
   19316: out<=1;
   19317: out<=1;
   19318: out<=1;
   19319: out<=1;
   19320: out<=1;
   19321: out<=1;
   19322: out<=0;
   19323: out<=0;
   19324: out<=0;
   19325: out<=1;
   19326: out<=0;
   19327: out<=1;
   19328: out<=1;
   19329: out<=0;
   19330: out<=0;
   19331: out<=1;
   19332: out<=0;
   19333: out<=0;
   19334: out<=0;
   19335: out<=0;
   19336: out<=0;
   19337: out<=0;
   19338: out<=1;
   19339: out<=1;
   19340: out<=1;
   19341: out<=0;
   19342: out<=1;
   19343: out<=0;
   19344: out<=0;
   19345: out<=1;
   19346: out<=1;
   19347: out<=0;
   19348: out<=1;
   19349: out<=1;
   19350: out<=1;
   19351: out<=1;
   19352: out<=1;
   19353: out<=1;
   19354: out<=0;
   19355: out<=0;
   19356: out<=0;
   19357: out<=1;
   19358: out<=0;
   19359: out<=1;
   19360: out<=1;
   19361: out<=0;
   19362: out<=0;
   19363: out<=1;
   19364: out<=0;
   19365: out<=0;
   19366: out<=0;
   19367: out<=0;
   19368: out<=0;
   19369: out<=0;
   19370: out<=1;
   19371: out<=1;
   19372: out<=1;
   19373: out<=0;
   19374: out<=1;
   19375: out<=0;
   19376: out<=0;
   19377: out<=1;
   19378: out<=1;
   19379: out<=0;
   19380: out<=1;
   19381: out<=1;
   19382: out<=1;
   19383: out<=1;
   19384: out<=1;
   19385: out<=1;
   19386: out<=0;
   19387: out<=0;
   19388: out<=0;
   19389: out<=1;
   19390: out<=0;
   19391: out<=1;
   19392: out<=0;
   19393: out<=1;
   19394: out<=1;
   19395: out<=0;
   19396: out<=1;
   19397: out<=1;
   19398: out<=1;
   19399: out<=1;
   19400: out<=1;
   19401: out<=1;
   19402: out<=0;
   19403: out<=0;
   19404: out<=0;
   19405: out<=1;
   19406: out<=0;
   19407: out<=1;
   19408: out<=0;
   19409: out<=1;
   19410: out<=1;
   19411: out<=0;
   19412: out<=1;
   19413: out<=1;
   19414: out<=1;
   19415: out<=1;
   19416: out<=1;
   19417: out<=1;
   19418: out<=0;
   19419: out<=0;
   19420: out<=0;
   19421: out<=1;
   19422: out<=0;
   19423: out<=1;
   19424: out<=1;
   19425: out<=0;
   19426: out<=0;
   19427: out<=1;
   19428: out<=0;
   19429: out<=0;
   19430: out<=0;
   19431: out<=0;
   19432: out<=0;
   19433: out<=0;
   19434: out<=1;
   19435: out<=1;
   19436: out<=1;
   19437: out<=0;
   19438: out<=1;
   19439: out<=0;
   19440: out<=1;
   19441: out<=0;
   19442: out<=0;
   19443: out<=1;
   19444: out<=0;
   19445: out<=0;
   19446: out<=0;
   19447: out<=0;
   19448: out<=0;
   19449: out<=0;
   19450: out<=1;
   19451: out<=1;
   19452: out<=1;
   19453: out<=0;
   19454: out<=1;
   19455: out<=0;
   19456: out<=0;
   19457: out<=0;
   19458: out<=1;
   19459: out<=1;
   19460: out<=1;
   19461: out<=0;
   19462: out<=1;
   19463: out<=0;
   19464: out<=0;
   19465: out<=1;
   19466: out<=1;
   19467: out<=0;
   19468: out<=1;
   19469: out<=1;
   19470: out<=1;
   19471: out<=1;
   19472: out<=0;
   19473: out<=0;
   19474: out<=1;
   19475: out<=1;
   19476: out<=1;
   19477: out<=0;
   19478: out<=1;
   19479: out<=0;
   19480: out<=0;
   19481: out<=1;
   19482: out<=1;
   19483: out<=0;
   19484: out<=1;
   19485: out<=1;
   19486: out<=1;
   19487: out<=1;
   19488: out<=1;
   19489: out<=1;
   19490: out<=0;
   19491: out<=0;
   19492: out<=0;
   19493: out<=1;
   19494: out<=0;
   19495: out<=1;
   19496: out<=1;
   19497: out<=0;
   19498: out<=0;
   19499: out<=1;
   19500: out<=0;
   19501: out<=0;
   19502: out<=0;
   19503: out<=0;
   19504: out<=1;
   19505: out<=1;
   19506: out<=0;
   19507: out<=0;
   19508: out<=0;
   19509: out<=1;
   19510: out<=0;
   19511: out<=1;
   19512: out<=1;
   19513: out<=0;
   19514: out<=0;
   19515: out<=1;
   19516: out<=0;
   19517: out<=0;
   19518: out<=0;
   19519: out<=0;
   19520: out<=1;
   19521: out<=1;
   19522: out<=0;
   19523: out<=0;
   19524: out<=0;
   19525: out<=1;
   19526: out<=0;
   19527: out<=1;
   19528: out<=1;
   19529: out<=0;
   19530: out<=0;
   19531: out<=1;
   19532: out<=0;
   19533: out<=0;
   19534: out<=0;
   19535: out<=0;
   19536: out<=0;
   19537: out<=0;
   19538: out<=1;
   19539: out<=1;
   19540: out<=1;
   19541: out<=0;
   19542: out<=1;
   19543: out<=0;
   19544: out<=0;
   19545: out<=1;
   19546: out<=1;
   19547: out<=0;
   19548: out<=1;
   19549: out<=1;
   19550: out<=1;
   19551: out<=1;
   19552: out<=1;
   19553: out<=1;
   19554: out<=0;
   19555: out<=0;
   19556: out<=0;
   19557: out<=1;
   19558: out<=0;
   19559: out<=1;
   19560: out<=1;
   19561: out<=0;
   19562: out<=0;
   19563: out<=1;
   19564: out<=0;
   19565: out<=0;
   19566: out<=0;
   19567: out<=0;
   19568: out<=0;
   19569: out<=0;
   19570: out<=1;
   19571: out<=1;
   19572: out<=1;
   19573: out<=0;
   19574: out<=1;
   19575: out<=0;
   19576: out<=0;
   19577: out<=1;
   19578: out<=1;
   19579: out<=0;
   19580: out<=1;
   19581: out<=1;
   19582: out<=1;
   19583: out<=1;
   19584: out<=0;
   19585: out<=0;
   19586: out<=1;
   19587: out<=1;
   19588: out<=1;
   19589: out<=0;
   19590: out<=1;
   19591: out<=0;
   19592: out<=0;
   19593: out<=1;
   19594: out<=1;
   19595: out<=0;
   19596: out<=1;
   19597: out<=1;
   19598: out<=1;
   19599: out<=1;
   19600: out<=1;
   19601: out<=1;
   19602: out<=0;
   19603: out<=0;
   19604: out<=0;
   19605: out<=1;
   19606: out<=0;
   19607: out<=1;
   19608: out<=1;
   19609: out<=0;
   19610: out<=0;
   19611: out<=1;
   19612: out<=0;
   19613: out<=0;
   19614: out<=0;
   19615: out<=0;
   19616: out<=1;
   19617: out<=1;
   19618: out<=0;
   19619: out<=0;
   19620: out<=0;
   19621: out<=1;
   19622: out<=0;
   19623: out<=1;
   19624: out<=1;
   19625: out<=0;
   19626: out<=0;
   19627: out<=1;
   19628: out<=0;
   19629: out<=0;
   19630: out<=0;
   19631: out<=0;
   19632: out<=0;
   19633: out<=0;
   19634: out<=1;
   19635: out<=1;
   19636: out<=1;
   19637: out<=0;
   19638: out<=1;
   19639: out<=0;
   19640: out<=0;
   19641: out<=1;
   19642: out<=1;
   19643: out<=0;
   19644: out<=1;
   19645: out<=1;
   19646: out<=1;
   19647: out<=1;
   19648: out<=1;
   19649: out<=1;
   19650: out<=0;
   19651: out<=0;
   19652: out<=0;
   19653: out<=1;
   19654: out<=0;
   19655: out<=1;
   19656: out<=1;
   19657: out<=0;
   19658: out<=0;
   19659: out<=1;
   19660: out<=0;
   19661: out<=0;
   19662: out<=0;
   19663: out<=0;
   19664: out<=1;
   19665: out<=1;
   19666: out<=0;
   19667: out<=0;
   19668: out<=0;
   19669: out<=1;
   19670: out<=0;
   19671: out<=1;
   19672: out<=1;
   19673: out<=0;
   19674: out<=0;
   19675: out<=1;
   19676: out<=0;
   19677: out<=0;
   19678: out<=0;
   19679: out<=0;
   19680: out<=1;
   19681: out<=1;
   19682: out<=0;
   19683: out<=0;
   19684: out<=0;
   19685: out<=1;
   19686: out<=0;
   19687: out<=1;
   19688: out<=1;
   19689: out<=0;
   19690: out<=0;
   19691: out<=1;
   19692: out<=0;
   19693: out<=0;
   19694: out<=0;
   19695: out<=0;
   19696: out<=1;
   19697: out<=1;
   19698: out<=0;
   19699: out<=0;
   19700: out<=0;
   19701: out<=1;
   19702: out<=0;
   19703: out<=1;
   19704: out<=1;
   19705: out<=0;
   19706: out<=0;
   19707: out<=1;
   19708: out<=0;
   19709: out<=0;
   19710: out<=0;
   19711: out<=0;
   19712: out<=0;
   19713: out<=1;
   19714: out<=0;
   19715: out<=1;
   19716: out<=0;
   19717: out<=0;
   19718: out<=1;
   19719: out<=1;
   19720: out<=1;
   19721: out<=1;
   19722: out<=1;
   19723: out<=1;
   19724: out<=1;
   19725: out<=0;
   19726: out<=0;
   19727: out<=1;
   19728: out<=1;
   19729: out<=0;
   19730: out<=1;
   19731: out<=0;
   19732: out<=1;
   19733: out<=1;
   19734: out<=0;
   19735: out<=0;
   19736: out<=0;
   19737: out<=0;
   19738: out<=0;
   19739: out<=0;
   19740: out<=0;
   19741: out<=1;
   19742: out<=1;
   19743: out<=0;
   19744: out<=0;
   19745: out<=1;
   19746: out<=0;
   19747: out<=1;
   19748: out<=0;
   19749: out<=0;
   19750: out<=1;
   19751: out<=1;
   19752: out<=1;
   19753: out<=1;
   19754: out<=1;
   19755: out<=1;
   19756: out<=1;
   19757: out<=0;
   19758: out<=0;
   19759: out<=1;
   19760: out<=1;
   19761: out<=0;
   19762: out<=1;
   19763: out<=0;
   19764: out<=1;
   19765: out<=1;
   19766: out<=0;
   19767: out<=0;
   19768: out<=0;
   19769: out<=0;
   19770: out<=0;
   19771: out<=0;
   19772: out<=0;
   19773: out<=1;
   19774: out<=1;
   19775: out<=0;
   19776: out<=1;
   19777: out<=0;
   19778: out<=1;
   19779: out<=0;
   19780: out<=1;
   19781: out<=1;
   19782: out<=0;
   19783: out<=0;
   19784: out<=0;
   19785: out<=0;
   19786: out<=0;
   19787: out<=0;
   19788: out<=0;
   19789: out<=1;
   19790: out<=1;
   19791: out<=0;
   19792: out<=1;
   19793: out<=0;
   19794: out<=1;
   19795: out<=0;
   19796: out<=1;
   19797: out<=1;
   19798: out<=0;
   19799: out<=0;
   19800: out<=0;
   19801: out<=0;
   19802: out<=0;
   19803: out<=0;
   19804: out<=0;
   19805: out<=1;
   19806: out<=1;
   19807: out<=0;
   19808: out<=0;
   19809: out<=1;
   19810: out<=0;
   19811: out<=1;
   19812: out<=0;
   19813: out<=0;
   19814: out<=1;
   19815: out<=1;
   19816: out<=1;
   19817: out<=1;
   19818: out<=1;
   19819: out<=1;
   19820: out<=1;
   19821: out<=0;
   19822: out<=0;
   19823: out<=1;
   19824: out<=0;
   19825: out<=1;
   19826: out<=0;
   19827: out<=1;
   19828: out<=0;
   19829: out<=0;
   19830: out<=1;
   19831: out<=1;
   19832: out<=1;
   19833: out<=1;
   19834: out<=1;
   19835: out<=1;
   19836: out<=1;
   19837: out<=0;
   19838: out<=0;
   19839: out<=1;
   19840: out<=0;
   19841: out<=1;
   19842: out<=0;
   19843: out<=1;
   19844: out<=0;
   19845: out<=0;
   19846: out<=1;
   19847: out<=1;
   19848: out<=1;
   19849: out<=1;
   19850: out<=1;
   19851: out<=1;
   19852: out<=1;
   19853: out<=0;
   19854: out<=0;
   19855: out<=1;
   19856: out<=0;
   19857: out<=1;
   19858: out<=0;
   19859: out<=1;
   19860: out<=0;
   19861: out<=0;
   19862: out<=1;
   19863: out<=1;
   19864: out<=1;
   19865: out<=1;
   19866: out<=1;
   19867: out<=1;
   19868: out<=1;
   19869: out<=0;
   19870: out<=0;
   19871: out<=1;
   19872: out<=0;
   19873: out<=1;
   19874: out<=0;
   19875: out<=1;
   19876: out<=0;
   19877: out<=0;
   19878: out<=1;
   19879: out<=1;
   19880: out<=1;
   19881: out<=1;
   19882: out<=1;
   19883: out<=1;
   19884: out<=1;
   19885: out<=0;
   19886: out<=0;
   19887: out<=1;
   19888: out<=0;
   19889: out<=1;
   19890: out<=0;
   19891: out<=1;
   19892: out<=0;
   19893: out<=0;
   19894: out<=1;
   19895: out<=1;
   19896: out<=1;
   19897: out<=1;
   19898: out<=1;
   19899: out<=1;
   19900: out<=1;
   19901: out<=0;
   19902: out<=0;
   19903: out<=1;
   19904: out<=1;
   19905: out<=0;
   19906: out<=1;
   19907: out<=0;
   19908: out<=1;
   19909: out<=1;
   19910: out<=0;
   19911: out<=0;
   19912: out<=0;
   19913: out<=0;
   19914: out<=0;
   19915: out<=0;
   19916: out<=0;
   19917: out<=1;
   19918: out<=1;
   19919: out<=0;
   19920: out<=0;
   19921: out<=1;
   19922: out<=0;
   19923: out<=1;
   19924: out<=0;
   19925: out<=0;
   19926: out<=1;
   19927: out<=1;
   19928: out<=1;
   19929: out<=1;
   19930: out<=1;
   19931: out<=1;
   19932: out<=1;
   19933: out<=0;
   19934: out<=0;
   19935: out<=1;
   19936: out<=0;
   19937: out<=1;
   19938: out<=0;
   19939: out<=1;
   19940: out<=0;
   19941: out<=0;
   19942: out<=1;
   19943: out<=1;
   19944: out<=1;
   19945: out<=1;
   19946: out<=1;
   19947: out<=1;
   19948: out<=1;
   19949: out<=0;
   19950: out<=0;
   19951: out<=1;
   19952: out<=1;
   19953: out<=0;
   19954: out<=1;
   19955: out<=0;
   19956: out<=1;
   19957: out<=1;
   19958: out<=0;
   19959: out<=0;
   19960: out<=0;
   19961: out<=0;
   19962: out<=0;
   19963: out<=0;
   19964: out<=0;
   19965: out<=1;
   19966: out<=1;
   19967: out<=0;
   19968: out<=1;
   19969: out<=0;
   19970: out<=0;
   19971: out<=1;
   19972: out<=1;
   19973: out<=1;
   19974: out<=1;
   19975: out<=1;
   19976: out<=1;
   19977: out<=1;
   19978: out<=0;
   19979: out<=0;
   19980: out<=1;
   19981: out<=0;
   19982: out<=1;
   19983: out<=0;
   19984: out<=0;
   19985: out<=1;
   19986: out<=1;
   19987: out<=0;
   19988: out<=0;
   19989: out<=0;
   19990: out<=0;
   19991: out<=0;
   19992: out<=0;
   19993: out<=0;
   19994: out<=1;
   19995: out<=1;
   19996: out<=0;
   19997: out<=1;
   19998: out<=0;
   19999: out<=1;
   20000: out<=0;
   20001: out<=1;
   20002: out<=1;
   20003: out<=0;
   20004: out<=0;
   20005: out<=0;
   20006: out<=0;
   20007: out<=0;
   20008: out<=0;
   20009: out<=0;
   20010: out<=1;
   20011: out<=1;
   20012: out<=0;
   20013: out<=1;
   20014: out<=0;
   20015: out<=1;
   20016: out<=1;
   20017: out<=0;
   20018: out<=0;
   20019: out<=1;
   20020: out<=1;
   20021: out<=1;
   20022: out<=1;
   20023: out<=1;
   20024: out<=1;
   20025: out<=1;
   20026: out<=0;
   20027: out<=0;
   20028: out<=1;
   20029: out<=0;
   20030: out<=1;
   20031: out<=0;
   20032: out<=0;
   20033: out<=1;
   20034: out<=1;
   20035: out<=0;
   20036: out<=0;
   20037: out<=0;
   20038: out<=0;
   20039: out<=0;
   20040: out<=0;
   20041: out<=0;
   20042: out<=1;
   20043: out<=1;
   20044: out<=0;
   20045: out<=1;
   20046: out<=0;
   20047: out<=1;
   20048: out<=0;
   20049: out<=1;
   20050: out<=1;
   20051: out<=0;
   20052: out<=0;
   20053: out<=0;
   20054: out<=0;
   20055: out<=0;
   20056: out<=0;
   20057: out<=0;
   20058: out<=1;
   20059: out<=1;
   20060: out<=0;
   20061: out<=1;
   20062: out<=0;
   20063: out<=1;
   20064: out<=0;
   20065: out<=1;
   20066: out<=1;
   20067: out<=0;
   20068: out<=0;
   20069: out<=0;
   20070: out<=0;
   20071: out<=0;
   20072: out<=0;
   20073: out<=0;
   20074: out<=1;
   20075: out<=1;
   20076: out<=0;
   20077: out<=1;
   20078: out<=0;
   20079: out<=1;
   20080: out<=0;
   20081: out<=1;
   20082: out<=1;
   20083: out<=0;
   20084: out<=0;
   20085: out<=0;
   20086: out<=0;
   20087: out<=0;
   20088: out<=0;
   20089: out<=0;
   20090: out<=1;
   20091: out<=1;
   20092: out<=0;
   20093: out<=1;
   20094: out<=0;
   20095: out<=1;
   20096: out<=1;
   20097: out<=0;
   20098: out<=0;
   20099: out<=1;
   20100: out<=1;
   20101: out<=1;
   20102: out<=1;
   20103: out<=1;
   20104: out<=1;
   20105: out<=1;
   20106: out<=0;
   20107: out<=0;
   20108: out<=1;
   20109: out<=0;
   20110: out<=1;
   20111: out<=0;
   20112: out<=1;
   20113: out<=0;
   20114: out<=0;
   20115: out<=1;
   20116: out<=1;
   20117: out<=1;
   20118: out<=1;
   20119: out<=1;
   20120: out<=1;
   20121: out<=1;
   20122: out<=0;
   20123: out<=0;
   20124: out<=1;
   20125: out<=0;
   20126: out<=1;
   20127: out<=0;
   20128: out<=0;
   20129: out<=1;
   20130: out<=1;
   20131: out<=0;
   20132: out<=0;
   20133: out<=0;
   20134: out<=0;
   20135: out<=0;
   20136: out<=0;
   20137: out<=0;
   20138: out<=1;
   20139: out<=1;
   20140: out<=0;
   20141: out<=1;
   20142: out<=0;
   20143: out<=1;
   20144: out<=0;
   20145: out<=1;
   20146: out<=1;
   20147: out<=0;
   20148: out<=0;
   20149: out<=0;
   20150: out<=0;
   20151: out<=0;
   20152: out<=0;
   20153: out<=0;
   20154: out<=1;
   20155: out<=1;
   20156: out<=0;
   20157: out<=1;
   20158: out<=0;
   20159: out<=1;
   20160: out<=0;
   20161: out<=1;
   20162: out<=1;
   20163: out<=0;
   20164: out<=0;
   20165: out<=0;
   20166: out<=0;
   20167: out<=0;
   20168: out<=0;
   20169: out<=0;
   20170: out<=1;
   20171: out<=1;
   20172: out<=0;
   20173: out<=1;
   20174: out<=0;
   20175: out<=1;
   20176: out<=1;
   20177: out<=0;
   20178: out<=0;
   20179: out<=1;
   20180: out<=1;
   20181: out<=1;
   20182: out<=1;
   20183: out<=1;
   20184: out<=1;
   20185: out<=1;
   20186: out<=0;
   20187: out<=0;
   20188: out<=1;
   20189: out<=0;
   20190: out<=1;
   20191: out<=0;
   20192: out<=0;
   20193: out<=1;
   20194: out<=1;
   20195: out<=0;
   20196: out<=0;
   20197: out<=0;
   20198: out<=0;
   20199: out<=0;
   20200: out<=0;
   20201: out<=0;
   20202: out<=1;
   20203: out<=1;
   20204: out<=0;
   20205: out<=1;
   20206: out<=0;
   20207: out<=1;
   20208: out<=1;
   20209: out<=0;
   20210: out<=0;
   20211: out<=1;
   20212: out<=1;
   20213: out<=1;
   20214: out<=1;
   20215: out<=1;
   20216: out<=1;
   20217: out<=1;
   20218: out<=0;
   20219: out<=0;
   20220: out<=1;
   20221: out<=0;
   20222: out<=1;
   20223: out<=0;
   20224: out<=1;
   20225: out<=1;
   20226: out<=1;
   20227: out<=1;
   20228: out<=0;
   20229: out<=1;
   20230: out<=1;
   20231: out<=0;
   20232: out<=0;
   20233: out<=1;
   20234: out<=0;
   20235: out<=1;
   20236: out<=1;
   20237: out<=1;
   20238: out<=0;
   20239: out<=0;
   20240: out<=1;
   20241: out<=1;
   20242: out<=1;
   20243: out<=1;
   20244: out<=0;
   20245: out<=1;
   20246: out<=1;
   20247: out<=0;
   20248: out<=0;
   20249: out<=1;
   20250: out<=0;
   20251: out<=1;
   20252: out<=1;
   20253: out<=1;
   20254: out<=0;
   20255: out<=0;
   20256: out<=1;
   20257: out<=1;
   20258: out<=1;
   20259: out<=1;
   20260: out<=0;
   20261: out<=1;
   20262: out<=1;
   20263: out<=0;
   20264: out<=0;
   20265: out<=1;
   20266: out<=0;
   20267: out<=1;
   20268: out<=1;
   20269: out<=1;
   20270: out<=0;
   20271: out<=0;
   20272: out<=1;
   20273: out<=1;
   20274: out<=1;
   20275: out<=1;
   20276: out<=0;
   20277: out<=1;
   20278: out<=1;
   20279: out<=0;
   20280: out<=0;
   20281: out<=1;
   20282: out<=0;
   20283: out<=1;
   20284: out<=1;
   20285: out<=1;
   20286: out<=0;
   20287: out<=0;
   20288: out<=0;
   20289: out<=0;
   20290: out<=0;
   20291: out<=0;
   20292: out<=1;
   20293: out<=0;
   20294: out<=0;
   20295: out<=1;
   20296: out<=1;
   20297: out<=0;
   20298: out<=1;
   20299: out<=0;
   20300: out<=0;
   20301: out<=0;
   20302: out<=1;
   20303: out<=1;
   20304: out<=1;
   20305: out<=1;
   20306: out<=1;
   20307: out<=1;
   20308: out<=0;
   20309: out<=1;
   20310: out<=1;
   20311: out<=0;
   20312: out<=0;
   20313: out<=1;
   20314: out<=0;
   20315: out<=1;
   20316: out<=1;
   20317: out<=1;
   20318: out<=0;
   20319: out<=0;
   20320: out<=1;
   20321: out<=1;
   20322: out<=1;
   20323: out<=1;
   20324: out<=0;
   20325: out<=1;
   20326: out<=1;
   20327: out<=0;
   20328: out<=0;
   20329: out<=1;
   20330: out<=0;
   20331: out<=1;
   20332: out<=1;
   20333: out<=1;
   20334: out<=0;
   20335: out<=0;
   20336: out<=0;
   20337: out<=0;
   20338: out<=0;
   20339: out<=0;
   20340: out<=1;
   20341: out<=0;
   20342: out<=0;
   20343: out<=1;
   20344: out<=1;
   20345: out<=0;
   20346: out<=1;
   20347: out<=0;
   20348: out<=0;
   20349: out<=0;
   20350: out<=1;
   20351: out<=1;
   20352: out<=1;
   20353: out<=1;
   20354: out<=1;
   20355: out<=1;
   20356: out<=0;
   20357: out<=1;
   20358: out<=1;
   20359: out<=0;
   20360: out<=0;
   20361: out<=1;
   20362: out<=0;
   20363: out<=1;
   20364: out<=1;
   20365: out<=1;
   20366: out<=0;
   20367: out<=0;
   20368: out<=0;
   20369: out<=0;
   20370: out<=0;
   20371: out<=0;
   20372: out<=1;
   20373: out<=0;
   20374: out<=0;
   20375: out<=1;
   20376: out<=1;
   20377: out<=0;
   20378: out<=1;
   20379: out<=0;
   20380: out<=0;
   20381: out<=0;
   20382: out<=1;
   20383: out<=1;
   20384: out<=1;
   20385: out<=1;
   20386: out<=1;
   20387: out<=1;
   20388: out<=0;
   20389: out<=1;
   20390: out<=1;
   20391: out<=0;
   20392: out<=0;
   20393: out<=1;
   20394: out<=0;
   20395: out<=1;
   20396: out<=1;
   20397: out<=1;
   20398: out<=0;
   20399: out<=0;
   20400: out<=0;
   20401: out<=0;
   20402: out<=0;
   20403: out<=0;
   20404: out<=1;
   20405: out<=0;
   20406: out<=0;
   20407: out<=1;
   20408: out<=1;
   20409: out<=0;
   20410: out<=1;
   20411: out<=0;
   20412: out<=0;
   20413: out<=0;
   20414: out<=1;
   20415: out<=1;
   20416: out<=0;
   20417: out<=0;
   20418: out<=0;
   20419: out<=0;
   20420: out<=1;
   20421: out<=0;
   20422: out<=0;
   20423: out<=1;
   20424: out<=1;
   20425: out<=0;
   20426: out<=1;
   20427: out<=0;
   20428: out<=0;
   20429: out<=0;
   20430: out<=1;
   20431: out<=1;
   20432: out<=0;
   20433: out<=0;
   20434: out<=0;
   20435: out<=0;
   20436: out<=1;
   20437: out<=0;
   20438: out<=0;
   20439: out<=1;
   20440: out<=1;
   20441: out<=0;
   20442: out<=1;
   20443: out<=0;
   20444: out<=0;
   20445: out<=0;
   20446: out<=1;
   20447: out<=1;
   20448: out<=1;
   20449: out<=1;
   20450: out<=1;
   20451: out<=1;
   20452: out<=0;
   20453: out<=1;
   20454: out<=1;
   20455: out<=0;
   20456: out<=0;
   20457: out<=1;
   20458: out<=0;
   20459: out<=1;
   20460: out<=1;
   20461: out<=1;
   20462: out<=0;
   20463: out<=0;
   20464: out<=1;
   20465: out<=1;
   20466: out<=1;
   20467: out<=1;
   20468: out<=0;
   20469: out<=1;
   20470: out<=1;
   20471: out<=0;
   20472: out<=0;
   20473: out<=1;
   20474: out<=0;
   20475: out<=1;
   20476: out<=1;
   20477: out<=1;
   20478: out<=0;
   20479: out<=0;
   20480: out<=1;
   20481: out<=0;
   20482: out<=0;
   20483: out<=1;
   20484: out<=0;
   20485: out<=0;
   20486: out<=0;
   20487: out<=0;
   20488: out<=1;
   20489: out<=1;
   20490: out<=0;
   20491: out<=0;
   20492: out<=0;
   20493: out<=1;
   20494: out<=0;
   20495: out<=1;
   20496: out<=0;
   20497: out<=1;
   20498: out<=1;
   20499: out<=0;
   20500: out<=1;
   20501: out<=1;
   20502: out<=1;
   20503: out<=1;
   20504: out<=0;
   20505: out<=0;
   20506: out<=1;
   20507: out<=1;
   20508: out<=1;
   20509: out<=0;
   20510: out<=1;
   20511: out<=0;
   20512: out<=1;
   20513: out<=0;
   20514: out<=0;
   20515: out<=1;
   20516: out<=0;
   20517: out<=0;
   20518: out<=0;
   20519: out<=0;
   20520: out<=1;
   20521: out<=1;
   20522: out<=0;
   20523: out<=0;
   20524: out<=0;
   20525: out<=1;
   20526: out<=0;
   20527: out<=1;
   20528: out<=0;
   20529: out<=1;
   20530: out<=1;
   20531: out<=0;
   20532: out<=1;
   20533: out<=1;
   20534: out<=1;
   20535: out<=1;
   20536: out<=0;
   20537: out<=0;
   20538: out<=1;
   20539: out<=1;
   20540: out<=1;
   20541: out<=0;
   20542: out<=1;
   20543: out<=0;
   20544: out<=1;
   20545: out<=0;
   20546: out<=0;
   20547: out<=1;
   20548: out<=0;
   20549: out<=0;
   20550: out<=0;
   20551: out<=0;
   20552: out<=1;
   20553: out<=1;
   20554: out<=0;
   20555: out<=0;
   20556: out<=0;
   20557: out<=1;
   20558: out<=0;
   20559: out<=1;
   20560: out<=1;
   20561: out<=0;
   20562: out<=0;
   20563: out<=1;
   20564: out<=0;
   20565: out<=0;
   20566: out<=0;
   20567: out<=0;
   20568: out<=1;
   20569: out<=1;
   20570: out<=0;
   20571: out<=0;
   20572: out<=0;
   20573: out<=1;
   20574: out<=0;
   20575: out<=1;
   20576: out<=0;
   20577: out<=1;
   20578: out<=1;
   20579: out<=0;
   20580: out<=1;
   20581: out<=1;
   20582: out<=1;
   20583: out<=1;
   20584: out<=0;
   20585: out<=0;
   20586: out<=1;
   20587: out<=1;
   20588: out<=1;
   20589: out<=0;
   20590: out<=1;
   20591: out<=0;
   20592: out<=0;
   20593: out<=1;
   20594: out<=1;
   20595: out<=0;
   20596: out<=1;
   20597: out<=1;
   20598: out<=1;
   20599: out<=1;
   20600: out<=0;
   20601: out<=0;
   20602: out<=1;
   20603: out<=1;
   20604: out<=1;
   20605: out<=0;
   20606: out<=1;
   20607: out<=0;
   20608: out<=0;
   20609: out<=1;
   20610: out<=1;
   20611: out<=0;
   20612: out<=1;
   20613: out<=1;
   20614: out<=1;
   20615: out<=1;
   20616: out<=0;
   20617: out<=0;
   20618: out<=1;
   20619: out<=1;
   20620: out<=1;
   20621: out<=0;
   20622: out<=1;
   20623: out<=0;
   20624: out<=0;
   20625: out<=1;
   20626: out<=1;
   20627: out<=0;
   20628: out<=1;
   20629: out<=1;
   20630: out<=1;
   20631: out<=1;
   20632: out<=0;
   20633: out<=0;
   20634: out<=1;
   20635: out<=1;
   20636: out<=1;
   20637: out<=0;
   20638: out<=1;
   20639: out<=0;
   20640: out<=0;
   20641: out<=1;
   20642: out<=1;
   20643: out<=0;
   20644: out<=1;
   20645: out<=1;
   20646: out<=1;
   20647: out<=1;
   20648: out<=0;
   20649: out<=0;
   20650: out<=1;
   20651: out<=1;
   20652: out<=1;
   20653: out<=0;
   20654: out<=1;
   20655: out<=0;
   20656: out<=0;
   20657: out<=1;
   20658: out<=1;
   20659: out<=0;
   20660: out<=1;
   20661: out<=1;
   20662: out<=1;
   20663: out<=1;
   20664: out<=0;
   20665: out<=0;
   20666: out<=1;
   20667: out<=1;
   20668: out<=1;
   20669: out<=0;
   20670: out<=1;
   20671: out<=0;
   20672: out<=0;
   20673: out<=1;
   20674: out<=1;
   20675: out<=0;
   20676: out<=1;
   20677: out<=1;
   20678: out<=1;
   20679: out<=1;
   20680: out<=0;
   20681: out<=0;
   20682: out<=1;
   20683: out<=1;
   20684: out<=1;
   20685: out<=0;
   20686: out<=1;
   20687: out<=0;
   20688: out<=1;
   20689: out<=0;
   20690: out<=0;
   20691: out<=1;
   20692: out<=0;
   20693: out<=0;
   20694: out<=0;
   20695: out<=0;
   20696: out<=1;
   20697: out<=1;
   20698: out<=0;
   20699: out<=0;
   20700: out<=0;
   20701: out<=1;
   20702: out<=0;
   20703: out<=1;
   20704: out<=1;
   20705: out<=0;
   20706: out<=0;
   20707: out<=1;
   20708: out<=0;
   20709: out<=0;
   20710: out<=0;
   20711: out<=0;
   20712: out<=1;
   20713: out<=1;
   20714: out<=0;
   20715: out<=0;
   20716: out<=0;
   20717: out<=1;
   20718: out<=0;
   20719: out<=1;
   20720: out<=0;
   20721: out<=1;
   20722: out<=1;
   20723: out<=0;
   20724: out<=1;
   20725: out<=1;
   20726: out<=1;
   20727: out<=1;
   20728: out<=0;
   20729: out<=0;
   20730: out<=1;
   20731: out<=1;
   20732: out<=1;
   20733: out<=0;
   20734: out<=1;
   20735: out<=0;
   20736: out<=1;
   20737: out<=1;
   20738: out<=1;
   20739: out<=1;
   20740: out<=1;
   20741: out<=0;
   20742: out<=0;
   20743: out<=1;
   20744: out<=0;
   20745: out<=1;
   20746: out<=0;
   20747: out<=1;
   20748: out<=0;
   20749: out<=0;
   20750: out<=1;
   20751: out<=1;
   20752: out<=1;
   20753: out<=1;
   20754: out<=1;
   20755: out<=1;
   20756: out<=1;
   20757: out<=0;
   20758: out<=0;
   20759: out<=1;
   20760: out<=0;
   20761: out<=1;
   20762: out<=0;
   20763: out<=1;
   20764: out<=0;
   20765: out<=0;
   20766: out<=1;
   20767: out<=1;
   20768: out<=0;
   20769: out<=0;
   20770: out<=0;
   20771: out<=0;
   20772: out<=0;
   20773: out<=1;
   20774: out<=1;
   20775: out<=0;
   20776: out<=1;
   20777: out<=0;
   20778: out<=1;
   20779: out<=0;
   20780: out<=1;
   20781: out<=1;
   20782: out<=0;
   20783: out<=0;
   20784: out<=0;
   20785: out<=0;
   20786: out<=0;
   20787: out<=0;
   20788: out<=0;
   20789: out<=1;
   20790: out<=1;
   20791: out<=0;
   20792: out<=1;
   20793: out<=0;
   20794: out<=1;
   20795: out<=0;
   20796: out<=1;
   20797: out<=1;
   20798: out<=0;
   20799: out<=0;
   20800: out<=1;
   20801: out<=1;
   20802: out<=1;
   20803: out<=1;
   20804: out<=1;
   20805: out<=0;
   20806: out<=0;
   20807: out<=1;
   20808: out<=0;
   20809: out<=1;
   20810: out<=0;
   20811: out<=1;
   20812: out<=0;
   20813: out<=0;
   20814: out<=1;
   20815: out<=1;
   20816: out<=0;
   20817: out<=0;
   20818: out<=0;
   20819: out<=0;
   20820: out<=0;
   20821: out<=1;
   20822: out<=1;
   20823: out<=0;
   20824: out<=1;
   20825: out<=0;
   20826: out<=1;
   20827: out<=0;
   20828: out<=1;
   20829: out<=1;
   20830: out<=0;
   20831: out<=0;
   20832: out<=1;
   20833: out<=1;
   20834: out<=1;
   20835: out<=1;
   20836: out<=1;
   20837: out<=0;
   20838: out<=0;
   20839: out<=1;
   20840: out<=0;
   20841: out<=1;
   20842: out<=0;
   20843: out<=1;
   20844: out<=0;
   20845: out<=0;
   20846: out<=1;
   20847: out<=1;
   20848: out<=0;
   20849: out<=0;
   20850: out<=0;
   20851: out<=0;
   20852: out<=0;
   20853: out<=1;
   20854: out<=1;
   20855: out<=0;
   20856: out<=1;
   20857: out<=0;
   20858: out<=1;
   20859: out<=0;
   20860: out<=1;
   20861: out<=1;
   20862: out<=0;
   20863: out<=0;
   20864: out<=0;
   20865: out<=0;
   20866: out<=0;
   20867: out<=0;
   20868: out<=0;
   20869: out<=1;
   20870: out<=1;
   20871: out<=0;
   20872: out<=1;
   20873: out<=0;
   20874: out<=1;
   20875: out<=0;
   20876: out<=1;
   20877: out<=1;
   20878: out<=0;
   20879: out<=0;
   20880: out<=1;
   20881: out<=1;
   20882: out<=1;
   20883: out<=1;
   20884: out<=1;
   20885: out<=0;
   20886: out<=0;
   20887: out<=1;
   20888: out<=0;
   20889: out<=1;
   20890: out<=0;
   20891: out<=1;
   20892: out<=0;
   20893: out<=0;
   20894: out<=1;
   20895: out<=1;
   20896: out<=1;
   20897: out<=1;
   20898: out<=1;
   20899: out<=1;
   20900: out<=1;
   20901: out<=0;
   20902: out<=0;
   20903: out<=1;
   20904: out<=0;
   20905: out<=1;
   20906: out<=0;
   20907: out<=1;
   20908: out<=0;
   20909: out<=0;
   20910: out<=1;
   20911: out<=1;
   20912: out<=0;
   20913: out<=0;
   20914: out<=0;
   20915: out<=0;
   20916: out<=0;
   20917: out<=1;
   20918: out<=1;
   20919: out<=0;
   20920: out<=1;
   20921: out<=0;
   20922: out<=1;
   20923: out<=0;
   20924: out<=1;
   20925: out<=1;
   20926: out<=0;
   20927: out<=0;
   20928: out<=0;
   20929: out<=0;
   20930: out<=0;
   20931: out<=0;
   20932: out<=0;
   20933: out<=1;
   20934: out<=1;
   20935: out<=0;
   20936: out<=1;
   20937: out<=0;
   20938: out<=1;
   20939: out<=0;
   20940: out<=1;
   20941: out<=1;
   20942: out<=0;
   20943: out<=0;
   20944: out<=0;
   20945: out<=0;
   20946: out<=0;
   20947: out<=0;
   20948: out<=0;
   20949: out<=1;
   20950: out<=1;
   20951: out<=0;
   20952: out<=1;
   20953: out<=0;
   20954: out<=1;
   20955: out<=0;
   20956: out<=1;
   20957: out<=1;
   20958: out<=0;
   20959: out<=0;
   20960: out<=0;
   20961: out<=0;
   20962: out<=0;
   20963: out<=0;
   20964: out<=0;
   20965: out<=1;
   20966: out<=1;
   20967: out<=0;
   20968: out<=1;
   20969: out<=0;
   20970: out<=1;
   20971: out<=0;
   20972: out<=1;
   20973: out<=1;
   20974: out<=0;
   20975: out<=0;
   20976: out<=0;
   20977: out<=0;
   20978: out<=0;
   20979: out<=0;
   20980: out<=0;
   20981: out<=1;
   20982: out<=1;
   20983: out<=0;
   20984: out<=1;
   20985: out<=0;
   20986: out<=1;
   20987: out<=0;
   20988: out<=1;
   20989: out<=1;
   20990: out<=0;
   20991: out<=0;
   20992: out<=1;
   20993: out<=1;
   20994: out<=0;
   20995: out<=0;
   20996: out<=1;
   20997: out<=0;
   20998: out<=1;
   20999: out<=0;
   21000: out<=1;
   21001: out<=0;
   21002: out<=0;
   21003: out<=1;
   21004: out<=1;
   21005: out<=1;
   21006: out<=1;
   21007: out<=1;
   21008: out<=1;
   21009: out<=1;
   21010: out<=0;
   21011: out<=0;
   21012: out<=1;
   21013: out<=0;
   21014: out<=1;
   21015: out<=0;
   21016: out<=1;
   21017: out<=0;
   21018: out<=0;
   21019: out<=1;
   21020: out<=1;
   21021: out<=1;
   21022: out<=1;
   21023: out<=1;
   21024: out<=1;
   21025: out<=1;
   21026: out<=0;
   21027: out<=0;
   21028: out<=1;
   21029: out<=0;
   21030: out<=1;
   21031: out<=0;
   21032: out<=1;
   21033: out<=0;
   21034: out<=0;
   21035: out<=1;
   21036: out<=1;
   21037: out<=1;
   21038: out<=1;
   21039: out<=1;
   21040: out<=1;
   21041: out<=1;
   21042: out<=0;
   21043: out<=0;
   21044: out<=1;
   21045: out<=0;
   21046: out<=1;
   21047: out<=0;
   21048: out<=1;
   21049: out<=0;
   21050: out<=0;
   21051: out<=1;
   21052: out<=1;
   21053: out<=1;
   21054: out<=1;
   21055: out<=1;
   21056: out<=1;
   21057: out<=1;
   21058: out<=0;
   21059: out<=0;
   21060: out<=1;
   21061: out<=0;
   21062: out<=1;
   21063: out<=0;
   21064: out<=1;
   21065: out<=0;
   21066: out<=0;
   21067: out<=1;
   21068: out<=1;
   21069: out<=1;
   21070: out<=1;
   21071: out<=1;
   21072: out<=0;
   21073: out<=0;
   21074: out<=1;
   21075: out<=1;
   21076: out<=0;
   21077: out<=1;
   21078: out<=0;
   21079: out<=1;
   21080: out<=0;
   21081: out<=1;
   21082: out<=1;
   21083: out<=0;
   21084: out<=0;
   21085: out<=0;
   21086: out<=0;
   21087: out<=0;
   21088: out<=0;
   21089: out<=0;
   21090: out<=1;
   21091: out<=1;
   21092: out<=0;
   21093: out<=1;
   21094: out<=0;
   21095: out<=1;
   21096: out<=0;
   21097: out<=1;
   21098: out<=1;
   21099: out<=0;
   21100: out<=0;
   21101: out<=0;
   21102: out<=0;
   21103: out<=0;
   21104: out<=1;
   21105: out<=1;
   21106: out<=0;
   21107: out<=0;
   21108: out<=1;
   21109: out<=0;
   21110: out<=1;
   21111: out<=0;
   21112: out<=1;
   21113: out<=0;
   21114: out<=0;
   21115: out<=1;
   21116: out<=1;
   21117: out<=1;
   21118: out<=1;
   21119: out<=1;
   21120: out<=0;
   21121: out<=0;
   21122: out<=1;
   21123: out<=1;
   21124: out<=0;
   21125: out<=1;
   21126: out<=0;
   21127: out<=1;
   21128: out<=0;
   21129: out<=1;
   21130: out<=1;
   21131: out<=0;
   21132: out<=0;
   21133: out<=0;
   21134: out<=0;
   21135: out<=0;
   21136: out<=1;
   21137: out<=1;
   21138: out<=0;
   21139: out<=0;
   21140: out<=1;
   21141: out<=0;
   21142: out<=1;
   21143: out<=0;
   21144: out<=1;
   21145: out<=0;
   21146: out<=0;
   21147: out<=1;
   21148: out<=1;
   21149: out<=1;
   21150: out<=1;
   21151: out<=1;
   21152: out<=0;
   21153: out<=0;
   21154: out<=1;
   21155: out<=1;
   21156: out<=0;
   21157: out<=1;
   21158: out<=0;
   21159: out<=1;
   21160: out<=0;
   21161: out<=1;
   21162: out<=1;
   21163: out<=0;
   21164: out<=0;
   21165: out<=0;
   21166: out<=0;
   21167: out<=0;
   21168: out<=1;
   21169: out<=1;
   21170: out<=0;
   21171: out<=0;
   21172: out<=1;
   21173: out<=0;
   21174: out<=1;
   21175: out<=0;
   21176: out<=1;
   21177: out<=0;
   21178: out<=0;
   21179: out<=1;
   21180: out<=1;
   21181: out<=1;
   21182: out<=1;
   21183: out<=1;
   21184: out<=0;
   21185: out<=0;
   21186: out<=1;
   21187: out<=1;
   21188: out<=0;
   21189: out<=1;
   21190: out<=0;
   21191: out<=1;
   21192: out<=0;
   21193: out<=1;
   21194: out<=1;
   21195: out<=0;
   21196: out<=0;
   21197: out<=0;
   21198: out<=0;
   21199: out<=0;
   21200: out<=0;
   21201: out<=0;
   21202: out<=1;
   21203: out<=1;
   21204: out<=0;
   21205: out<=1;
   21206: out<=0;
   21207: out<=1;
   21208: out<=0;
   21209: out<=1;
   21210: out<=1;
   21211: out<=0;
   21212: out<=0;
   21213: out<=0;
   21214: out<=0;
   21215: out<=0;
   21216: out<=1;
   21217: out<=1;
   21218: out<=0;
   21219: out<=0;
   21220: out<=1;
   21221: out<=0;
   21222: out<=1;
   21223: out<=0;
   21224: out<=1;
   21225: out<=0;
   21226: out<=0;
   21227: out<=1;
   21228: out<=1;
   21229: out<=1;
   21230: out<=1;
   21231: out<=1;
   21232: out<=1;
   21233: out<=1;
   21234: out<=0;
   21235: out<=0;
   21236: out<=1;
   21237: out<=0;
   21238: out<=1;
   21239: out<=0;
   21240: out<=1;
   21241: out<=0;
   21242: out<=0;
   21243: out<=1;
   21244: out<=1;
   21245: out<=1;
   21246: out<=1;
   21247: out<=1;
   21248: out<=1;
   21249: out<=0;
   21250: out<=1;
   21251: out<=0;
   21252: out<=0;
   21253: out<=0;
   21254: out<=1;
   21255: out<=1;
   21256: out<=0;
   21257: out<=0;
   21258: out<=0;
   21259: out<=0;
   21260: out<=1;
   21261: out<=0;
   21262: out<=0;
   21263: out<=1;
   21264: out<=0;
   21265: out<=1;
   21266: out<=0;
   21267: out<=1;
   21268: out<=1;
   21269: out<=1;
   21270: out<=0;
   21271: out<=0;
   21272: out<=1;
   21273: out<=1;
   21274: out<=1;
   21275: out<=1;
   21276: out<=0;
   21277: out<=1;
   21278: out<=1;
   21279: out<=0;
   21280: out<=0;
   21281: out<=1;
   21282: out<=0;
   21283: out<=1;
   21284: out<=1;
   21285: out<=1;
   21286: out<=0;
   21287: out<=0;
   21288: out<=1;
   21289: out<=1;
   21290: out<=1;
   21291: out<=1;
   21292: out<=0;
   21293: out<=1;
   21294: out<=1;
   21295: out<=0;
   21296: out<=1;
   21297: out<=0;
   21298: out<=1;
   21299: out<=0;
   21300: out<=0;
   21301: out<=0;
   21302: out<=1;
   21303: out<=1;
   21304: out<=0;
   21305: out<=0;
   21306: out<=0;
   21307: out<=0;
   21308: out<=1;
   21309: out<=0;
   21310: out<=0;
   21311: out<=1;
   21312: out<=1;
   21313: out<=0;
   21314: out<=1;
   21315: out<=0;
   21316: out<=0;
   21317: out<=0;
   21318: out<=1;
   21319: out<=1;
   21320: out<=0;
   21321: out<=0;
   21322: out<=0;
   21323: out<=0;
   21324: out<=1;
   21325: out<=0;
   21326: out<=0;
   21327: out<=1;
   21328: out<=1;
   21329: out<=0;
   21330: out<=1;
   21331: out<=0;
   21332: out<=0;
   21333: out<=0;
   21334: out<=1;
   21335: out<=1;
   21336: out<=0;
   21337: out<=0;
   21338: out<=0;
   21339: out<=0;
   21340: out<=1;
   21341: out<=0;
   21342: out<=0;
   21343: out<=1;
   21344: out<=1;
   21345: out<=0;
   21346: out<=1;
   21347: out<=0;
   21348: out<=0;
   21349: out<=0;
   21350: out<=1;
   21351: out<=1;
   21352: out<=0;
   21353: out<=0;
   21354: out<=0;
   21355: out<=0;
   21356: out<=1;
   21357: out<=0;
   21358: out<=0;
   21359: out<=1;
   21360: out<=1;
   21361: out<=0;
   21362: out<=1;
   21363: out<=0;
   21364: out<=0;
   21365: out<=0;
   21366: out<=1;
   21367: out<=1;
   21368: out<=0;
   21369: out<=0;
   21370: out<=0;
   21371: out<=0;
   21372: out<=1;
   21373: out<=0;
   21374: out<=0;
   21375: out<=1;
   21376: out<=0;
   21377: out<=1;
   21378: out<=0;
   21379: out<=1;
   21380: out<=1;
   21381: out<=1;
   21382: out<=0;
   21383: out<=0;
   21384: out<=1;
   21385: out<=1;
   21386: out<=1;
   21387: out<=1;
   21388: out<=0;
   21389: out<=1;
   21390: out<=1;
   21391: out<=0;
   21392: out<=0;
   21393: out<=1;
   21394: out<=0;
   21395: out<=1;
   21396: out<=1;
   21397: out<=1;
   21398: out<=0;
   21399: out<=0;
   21400: out<=1;
   21401: out<=1;
   21402: out<=1;
   21403: out<=1;
   21404: out<=0;
   21405: out<=1;
   21406: out<=1;
   21407: out<=0;
   21408: out<=1;
   21409: out<=0;
   21410: out<=1;
   21411: out<=0;
   21412: out<=0;
   21413: out<=0;
   21414: out<=1;
   21415: out<=1;
   21416: out<=0;
   21417: out<=0;
   21418: out<=0;
   21419: out<=0;
   21420: out<=1;
   21421: out<=0;
   21422: out<=0;
   21423: out<=1;
   21424: out<=1;
   21425: out<=0;
   21426: out<=1;
   21427: out<=0;
   21428: out<=0;
   21429: out<=0;
   21430: out<=1;
   21431: out<=1;
   21432: out<=0;
   21433: out<=0;
   21434: out<=0;
   21435: out<=0;
   21436: out<=1;
   21437: out<=0;
   21438: out<=0;
   21439: out<=1;
   21440: out<=0;
   21441: out<=1;
   21442: out<=0;
   21443: out<=1;
   21444: out<=1;
   21445: out<=1;
   21446: out<=0;
   21447: out<=0;
   21448: out<=1;
   21449: out<=1;
   21450: out<=1;
   21451: out<=1;
   21452: out<=0;
   21453: out<=1;
   21454: out<=1;
   21455: out<=0;
   21456: out<=1;
   21457: out<=0;
   21458: out<=1;
   21459: out<=0;
   21460: out<=0;
   21461: out<=0;
   21462: out<=1;
   21463: out<=1;
   21464: out<=0;
   21465: out<=0;
   21466: out<=0;
   21467: out<=0;
   21468: out<=1;
   21469: out<=0;
   21470: out<=0;
   21471: out<=1;
   21472: out<=0;
   21473: out<=1;
   21474: out<=0;
   21475: out<=1;
   21476: out<=1;
   21477: out<=1;
   21478: out<=0;
   21479: out<=0;
   21480: out<=1;
   21481: out<=1;
   21482: out<=1;
   21483: out<=1;
   21484: out<=0;
   21485: out<=1;
   21486: out<=1;
   21487: out<=0;
   21488: out<=1;
   21489: out<=0;
   21490: out<=1;
   21491: out<=0;
   21492: out<=0;
   21493: out<=0;
   21494: out<=1;
   21495: out<=1;
   21496: out<=0;
   21497: out<=0;
   21498: out<=0;
   21499: out<=0;
   21500: out<=1;
   21501: out<=0;
   21502: out<=0;
   21503: out<=1;
   21504: out<=1;
   21505: out<=1;
   21506: out<=1;
   21507: out<=1;
   21508: out<=0;
   21509: out<=1;
   21510: out<=1;
   21511: out<=0;
   21512: out<=1;
   21513: out<=0;
   21514: out<=1;
   21515: out<=0;
   21516: out<=0;
   21517: out<=0;
   21518: out<=1;
   21519: out<=1;
   21520: out<=0;
   21521: out<=0;
   21522: out<=0;
   21523: out<=0;
   21524: out<=1;
   21525: out<=0;
   21526: out<=0;
   21527: out<=1;
   21528: out<=0;
   21529: out<=1;
   21530: out<=0;
   21531: out<=1;
   21532: out<=1;
   21533: out<=1;
   21534: out<=0;
   21535: out<=0;
   21536: out<=1;
   21537: out<=1;
   21538: out<=1;
   21539: out<=1;
   21540: out<=0;
   21541: out<=1;
   21542: out<=1;
   21543: out<=0;
   21544: out<=1;
   21545: out<=0;
   21546: out<=1;
   21547: out<=0;
   21548: out<=0;
   21549: out<=0;
   21550: out<=1;
   21551: out<=1;
   21552: out<=0;
   21553: out<=0;
   21554: out<=0;
   21555: out<=0;
   21556: out<=1;
   21557: out<=0;
   21558: out<=0;
   21559: out<=1;
   21560: out<=0;
   21561: out<=1;
   21562: out<=0;
   21563: out<=1;
   21564: out<=1;
   21565: out<=1;
   21566: out<=0;
   21567: out<=0;
   21568: out<=1;
   21569: out<=1;
   21570: out<=1;
   21571: out<=1;
   21572: out<=0;
   21573: out<=1;
   21574: out<=1;
   21575: out<=0;
   21576: out<=1;
   21577: out<=0;
   21578: out<=1;
   21579: out<=0;
   21580: out<=0;
   21581: out<=0;
   21582: out<=1;
   21583: out<=1;
   21584: out<=1;
   21585: out<=1;
   21586: out<=1;
   21587: out<=1;
   21588: out<=0;
   21589: out<=1;
   21590: out<=1;
   21591: out<=0;
   21592: out<=1;
   21593: out<=0;
   21594: out<=1;
   21595: out<=0;
   21596: out<=0;
   21597: out<=0;
   21598: out<=1;
   21599: out<=1;
   21600: out<=0;
   21601: out<=0;
   21602: out<=0;
   21603: out<=0;
   21604: out<=1;
   21605: out<=0;
   21606: out<=0;
   21607: out<=1;
   21608: out<=0;
   21609: out<=1;
   21610: out<=0;
   21611: out<=1;
   21612: out<=1;
   21613: out<=1;
   21614: out<=0;
   21615: out<=0;
   21616: out<=0;
   21617: out<=0;
   21618: out<=0;
   21619: out<=0;
   21620: out<=1;
   21621: out<=0;
   21622: out<=0;
   21623: out<=1;
   21624: out<=0;
   21625: out<=1;
   21626: out<=0;
   21627: out<=1;
   21628: out<=1;
   21629: out<=1;
   21630: out<=0;
   21631: out<=0;
   21632: out<=0;
   21633: out<=0;
   21634: out<=0;
   21635: out<=0;
   21636: out<=1;
   21637: out<=0;
   21638: out<=0;
   21639: out<=1;
   21640: out<=0;
   21641: out<=1;
   21642: out<=0;
   21643: out<=1;
   21644: out<=1;
   21645: out<=1;
   21646: out<=0;
   21647: out<=0;
   21648: out<=0;
   21649: out<=0;
   21650: out<=0;
   21651: out<=0;
   21652: out<=1;
   21653: out<=0;
   21654: out<=0;
   21655: out<=1;
   21656: out<=0;
   21657: out<=1;
   21658: out<=0;
   21659: out<=1;
   21660: out<=1;
   21661: out<=1;
   21662: out<=0;
   21663: out<=0;
   21664: out<=0;
   21665: out<=0;
   21666: out<=0;
   21667: out<=0;
   21668: out<=1;
   21669: out<=0;
   21670: out<=0;
   21671: out<=1;
   21672: out<=0;
   21673: out<=1;
   21674: out<=0;
   21675: out<=1;
   21676: out<=1;
   21677: out<=1;
   21678: out<=0;
   21679: out<=0;
   21680: out<=0;
   21681: out<=0;
   21682: out<=0;
   21683: out<=0;
   21684: out<=1;
   21685: out<=0;
   21686: out<=0;
   21687: out<=1;
   21688: out<=0;
   21689: out<=1;
   21690: out<=0;
   21691: out<=1;
   21692: out<=1;
   21693: out<=1;
   21694: out<=0;
   21695: out<=0;
   21696: out<=0;
   21697: out<=0;
   21698: out<=0;
   21699: out<=0;
   21700: out<=1;
   21701: out<=0;
   21702: out<=0;
   21703: out<=1;
   21704: out<=0;
   21705: out<=1;
   21706: out<=0;
   21707: out<=1;
   21708: out<=1;
   21709: out<=1;
   21710: out<=0;
   21711: out<=0;
   21712: out<=1;
   21713: out<=1;
   21714: out<=1;
   21715: out<=1;
   21716: out<=0;
   21717: out<=1;
   21718: out<=1;
   21719: out<=0;
   21720: out<=1;
   21721: out<=0;
   21722: out<=1;
   21723: out<=0;
   21724: out<=0;
   21725: out<=0;
   21726: out<=1;
   21727: out<=1;
   21728: out<=1;
   21729: out<=1;
   21730: out<=1;
   21731: out<=1;
   21732: out<=0;
   21733: out<=1;
   21734: out<=1;
   21735: out<=0;
   21736: out<=1;
   21737: out<=0;
   21738: out<=1;
   21739: out<=0;
   21740: out<=0;
   21741: out<=0;
   21742: out<=1;
   21743: out<=1;
   21744: out<=0;
   21745: out<=0;
   21746: out<=0;
   21747: out<=0;
   21748: out<=1;
   21749: out<=0;
   21750: out<=0;
   21751: out<=1;
   21752: out<=0;
   21753: out<=1;
   21754: out<=0;
   21755: out<=1;
   21756: out<=1;
   21757: out<=1;
   21758: out<=0;
   21759: out<=0;
   21760: out<=0;
   21761: out<=1;
   21762: out<=1;
   21763: out<=0;
   21764: out<=0;
   21765: out<=0;
   21766: out<=0;
   21767: out<=0;
   21768: out<=1;
   21769: out<=1;
   21770: out<=0;
   21771: out<=0;
   21772: out<=1;
   21773: out<=0;
   21774: out<=1;
   21775: out<=0;
   21776: out<=0;
   21777: out<=1;
   21778: out<=1;
   21779: out<=0;
   21780: out<=0;
   21781: out<=0;
   21782: out<=0;
   21783: out<=0;
   21784: out<=1;
   21785: out<=1;
   21786: out<=0;
   21787: out<=0;
   21788: out<=1;
   21789: out<=0;
   21790: out<=1;
   21791: out<=0;
   21792: out<=1;
   21793: out<=0;
   21794: out<=0;
   21795: out<=1;
   21796: out<=1;
   21797: out<=1;
   21798: out<=1;
   21799: out<=1;
   21800: out<=0;
   21801: out<=0;
   21802: out<=1;
   21803: out<=1;
   21804: out<=0;
   21805: out<=1;
   21806: out<=0;
   21807: out<=1;
   21808: out<=1;
   21809: out<=0;
   21810: out<=0;
   21811: out<=1;
   21812: out<=1;
   21813: out<=1;
   21814: out<=1;
   21815: out<=1;
   21816: out<=0;
   21817: out<=0;
   21818: out<=1;
   21819: out<=1;
   21820: out<=0;
   21821: out<=1;
   21822: out<=0;
   21823: out<=1;
   21824: out<=0;
   21825: out<=1;
   21826: out<=1;
   21827: out<=0;
   21828: out<=0;
   21829: out<=0;
   21830: out<=0;
   21831: out<=0;
   21832: out<=1;
   21833: out<=1;
   21834: out<=0;
   21835: out<=0;
   21836: out<=1;
   21837: out<=0;
   21838: out<=1;
   21839: out<=0;
   21840: out<=1;
   21841: out<=0;
   21842: out<=0;
   21843: out<=1;
   21844: out<=1;
   21845: out<=1;
   21846: out<=1;
   21847: out<=1;
   21848: out<=0;
   21849: out<=0;
   21850: out<=1;
   21851: out<=1;
   21852: out<=0;
   21853: out<=1;
   21854: out<=0;
   21855: out<=1;
   21856: out<=0;
   21857: out<=1;
   21858: out<=1;
   21859: out<=0;
   21860: out<=0;
   21861: out<=0;
   21862: out<=0;
   21863: out<=0;
   21864: out<=1;
   21865: out<=1;
   21866: out<=0;
   21867: out<=0;
   21868: out<=1;
   21869: out<=0;
   21870: out<=1;
   21871: out<=0;
   21872: out<=1;
   21873: out<=0;
   21874: out<=0;
   21875: out<=1;
   21876: out<=1;
   21877: out<=1;
   21878: out<=1;
   21879: out<=1;
   21880: out<=0;
   21881: out<=0;
   21882: out<=1;
   21883: out<=1;
   21884: out<=0;
   21885: out<=1;
   21886: out<=0;
   21887: out<=1;
   21888: out<=1;
   21889: out<=0;
   21890: out<=0;
   21891: out<=1;
   21892: out<=1;
   21893: out<=1;
   21894: out<=1;
   21895: out<=1;
   21896: out<=0;
   21897: out<=0;
   21898: out<=1;
   21899: out<=1;
   21900: out<=0;
   21901: out<=1;
   21902: out<=0;
   21903: out<=1;
   21904: out<=0;
   21905: out<=1;
   21906: out<=1;
   21907: out<=0;
   21908: out<=0;
   21909: out<=0;
   21910: out<=0;
   21911: out<=0;
   21912: out<=1;
   21913: out<=1;
   21914: out<=0;
   21915: out<=0;
   21916: out<=1;
   21917: out<=0;
   21918: out<=1;
   21919: out<=0;
   21920: out<=0;
   21921: out<=1;
   21922: out<=1;
   21923: out<=0;
   21924: out<=0;
   21925: out<=0;
   21926: out<=0;
   21927: out<=0;
   21928: out<=1;
   21929: out<=1;
   21930: out<=0;
   21931: out<=0;
   21932: out<=1;
   21933: out<=0;
   21934: out<=1;
   21935: out<=0;
   21936: out<=1;
   21937: out<=0;
   21938: out<=0;
   21939: out<=1;
   21940: out<=1;
   21941: out<=1;
   21942: out<=1;
   21943: out<=1;
   21944: out<=0;
   21945: out<=0;
   21946: out<=1;
   21947: out<=1;
   21948: out<=0;
   21949: out<=1;
   21950: out<=0;
   21951: out<=1;
   21952: out<=1;
   21953: out<=0;
   21954: out<=0;
   21955: out<=1;
   21956: out<=1;
   21957: out<=1;
   21958: out<=1;
   21959: out<=1;
   21960: out<=0;
   21961: out<=0;
   21962: out<=1;
   21963: out<=1;
   21964: out<=0;
   21965: out<=1;
   21966: out<=0;
   21967: out<=1;
   21968: out<=1;
   21969: out<=0;
   21970: out<=0;
   21971: out<=1;
   21972: out<=1;
   21973: out<=1;
   21974: out<=1;
   21975: out<=1;
   21976: out<=0;
   21977: out<=0;
   21978: out<=1;
   21979: out<=1;
   21980: out<=0;
   21981: out<=1;
   21982: out<=0;
   21983: out<=1;
   21984: out<=1;
   21985: out<=0;
   21986: out<=0;
   21987: out<=1;
   21988: out<=1;
   21989: out<=1;
   21990: out<=1;
   21991: out<=1;
   21992: out<=0;
   21993: out<=0;
   21994: out<=1;
   21995: out<=1;
   21996: out<=0;
   21997: out<=1;
   21998: out<=0;
   21999: out<=1;
   22000: out<=1;
   22001: out<=0;
   22002: out<=0;
   22003: out<=1;
   22004: out<=1;
   22005: out<=1;
   22006: out<=1;
   22007: out<=1;
   22008: out<=0;
   22009: out<=0;
   22010: out<=1;
   22011: out<=1;
   22012: out<=0;
   22013: out<=1;
   22014: out<=0;
   22015: out<=1;
   22016: out<=0;
   22017: out<=1;
   22018: out<=0;
   22019: out<=1;
   22020: out<=0;
   22021: out<=0;
   22022: out<=1;
   22023: out<=1;
   22024: out<=0;
   22025: out<=0;
   22026: out<=0;
   22027: out<=0;
   22028: out<=0;
   22029: out<=1;
   22030: out<=1;
   22031: out<=0;
   22032: out<=0;
   22033: out<=1;
   22034: out<=0;
   22035: out<=1;
   22036: out<=0;
   22037: out<=0;
   22038: out<=1;
   22039: out<=1;
   22040: out<=0;
   22041: out<=0;
   22042: out<=0;
   22043: out<=0;
   22044: out<=0;
   22045: out<=1;
   22046: out<=1;
   22047: out<=0;
   22048: out<=0;
   22049: out<=1;
   22050: out<=0;
   22051: out<=1;
   22052: out<=0;
   22053: out<=0;
   22054: out<=1;
   22055: out<=1;
   22056: out<=0;
   22057: out<=0;
   22058: out<=0;
   22059: out<=0;
   22060: out<=0;
   22061: out<=1;
   22062: out<=1;
   22063: out<=0;
   22064: out<=0;
   22065: out<=1;
   22066: out<=0;
   22067: out<=1;
   22068: out<=0;
   22069: out<=0;
   22070: out<=1;
   22071: out<=1;
   22072: out<=0;
   22073: out<=0;
   22074: out<=0;
   22075: out<=0;
   22076: out<=0;
   22077: out<=1;
   22078: out<=1;
   22079: out<=0;
   22080: out<=0;
   22081: out<=1;
   22082: out<=0;
   22083: out<=1;
   22084: out<=0;
   22085: out<=0;
   22086: out<=1;
   22087: out<=1;
   22088: out<=0;
   22089: out<=0;
   22090: out<=0;
   22091: out<=0;
   22092: out<=0;
   22093: out<=1;
   22094: out<=1;
   22095: out<=0;
   22096: out<=1;
   22097: out<=0;
   22098: out<=1;
   22099: out<=0;
   22100: out<=1;
   22101: out<=1;
   22102: out<=0;
   22103: out<=0;
   22104: out<=1;
   22105: out<=1;
   22106: out<=1;
   22107: out<=1;
   22108: out<=1;
   22109: out<=0;
   22110: out<=0;
   22111: out<=1;
   22112: out<=1;
   22113: out<=0;
   22114: out<=1;
   22115: out<=0;
   22116: out<=1;
   22117: out<=1;
   22118: out<=0;
   22119: out<=0;
   22120: out<=1;
   22121: out<=1;
   22122: out<=1;
   22123: out<=1;
   22124: out<=1;
   22125: out<=0;
   22126: out<=0;
   22127: out<=1;
   22128: out<=0;
   22129: out<=1;
   22130: out<=0;
   22131: out<=1;
   22132: out<=0;
   22133: out<=0;
   22134: out<=1;
   22135: out<=1;
   22136: out<=0;
   22137: out<=0;
   22138: out<=0;
   22139: out<=0;
   22140: out<=0;
   22141: out<=1;
   22142: out<=1;
   22143: out<=0;
   22144: out<=1;
   22145: out<=0;
   22146: out<=1;
   22147: out<=0;
   22148: out<=1;
   22149: out<=1;
   22150: out<=0;
   22151: out<=0;
   22152: out<=1;
   22153: out<=1;
   22154: out<=1;
   22155: out<=1;
   22156: out<=1;
   22157: out<=0;
   22158: out<=0;
   22159: out<=1;
   22160: out<=0;
   22161: out<=1;
   22162: out<=0;
   22163: out<=1;
   22164: out<=0;
   22165: out<=0;
   22166: out<=1;
   22167: out<=1;
   22168: out<=0;
   22169: out<=0;
   22170: out<=0;
   22171: out<=0;
   22172: out<=0;
   22173: out<=1;
   22174: out<=1;
   22175: out<=0;
   22176: out<=1;
   22177: out<=0;
   22178: out<=1;
   22179: out<=0;
   22180: out<=1;
   22181: out<=1;
   22182: out<=0;
   22183: out<=0;
   22184: out<=1;
   22185: out<=1;
   22186: out<=1;
   22187: out<=1;
   22188: out<=1;
   22189: out<=0;
   22190: out<=0;
   22191: out<=1;
   22192: out<=0;
   22193: out<=1;
   22194: out<=0;
   22195: out<=1;
   22196: out<=0;
   22197: out<=0;
   22198: out<=1;
   22199: out<=1;
   22200: out<=0;
   22201: out<=0;
   22202: out<=0;
   22203: out<=0;
   22204: out<=0;
   22205: out<=1;
   22206: out<=1;
   22207: out<=0;
   22208: out<=1;
   22209: out<=0;
   22210: out<=1;
   22211: out<=0;
   22212: out<=1;
   22213: out<=1;
   22214: out<=0;
   22215: out<=0;
   22216: out<=1;
   22217: out<=1;
   22218: out<=1;
   22219: out<=1;
   22220: out<=1;
   22221: out<=0;
   22222: out<=0;
   22223: out<=1;
   22224: out<=1;
   22225: out<=0;
   22226: out<=1;
   22227: out<=0;
   22228: out<=1;
   22229: out<=1;
   22230: out<=0;
   22231: out<=0;
   22232: out<=1;
   22233: out<=1;
   22234: out<=1;
   22235: out<=1;
   22236: out<=1;
   22237: out<=0;
   22238: out<=0;
   22239: out<=1;
   22240: out<=0;
   22241: out<=1;
   22242: out<=0;
   22243: out<=1;
   22244: out<=0;
   22245: out<=0;
   22246: out<=1;
   22247: out<=1;
   22248: out<=0;
   22249: out<=0;
   22250: out<=0;
   22251: out<=0;
   22252: out<=0;
   22253: out<=1;
   22254: out<=1;
   22255: out<=0;
   22256: out<=0;
   22257: out<=1;
   22258: out<=0;
   22259: out<=1;
   22260: out<=0;
   22261: out<=0;
   22262: out<=1;
   22263: out<=1;
   22264: out<=0;
   22265: out<=0;
   22266: out<=0;
   22267: out<=0;
   22268: out<=0;
   22269: out<=1;
   22270: out<=1;
   22271: out<=0;
   22272: out<=1;
   22273: out<=1;
   22274: out<=0;
   22275: out<=0;
   22276: out<=0;
   22277: out<=1;
   22278: out<=0;
   22279: out<=1;
   22280: out<=0;
   22281: out<=1;
   22282: out<=1;
   22283: out<=0;
   22284: out<=1;
   22285: out<=1;
   22286: out<=1;
   22287: out<=1;
   22288: out<=0;
   22289: out<=0;
   22290: out<=1;
   22291: out<=1;
   22292: out<=1;
   22293: out<=0;
   22294: out<=1;
   22295: out<=0;
   22296: out<=1;
   22297: out<=0;
   22298: out<=0;
   22299: out<=1;
   22300: out<=0;
   22301: out<=0;
   22302: out<=0;
   22303: out<=0;
   22304: out<=0;
   22305: out<=0;
   22306: out<=1;
   22307: out<=1;
   22308: out<=1;
   22309: out<=0;
   22310: out<=1;
   22311: out<=0;
   22312: out<=1;
   22313: out<=0;
   22314: out<=0;
   22315: out<=1;
   22316: out<=0;
   22317: out<=0;
   22318: out<=0;
   22319: out<=0;
   22320: out<=1;
   22321: out<=1;
   22322: out<=0;
   22323: out<=0;
   22324: out<=0;
   22325: out<=1;
   22326: out<=0;
   22327: out<=1;
   22328: out<=0;
   22329: out<=1;
   22330: out<=1;
   22331: out<=0;
   22332: out<=1;
   22333: out<=1;
   22334: out<=1;
   22335: out<=1;
   22336: out<=1;
   22337: out<=1;
   22338: out<=0;
   22339: out<=0;
   22340: out<=0;
   22341: out<=1;
   22342: out<=0;
   22343: out<=1;
   22344: out<=0;
   22345: out<=1;
   22346: out<=1;
   22347: out<=0;
   22348: out<=1;
   22349: out<=1;
   22350: out<=1;
   22351: out<=1;
   22352: out<=1;
   22353: out<=1;
   22354: out<=0;
   22355: out<=0;
   22356: out<=0;
   22357: out<=1;
   22358: out<=0;
   22359: out<=1;
   22360: out<=0;
   22361: out<=1;
   22362: out<=1;
   22363: out<=0;
   22364: out<=1;
   22365: out<=1;
   22366: out<=1;
   22367: out<=1;
   22368: out<=1;
   22369: out<=1;
   22370: out<=0;
   22371: out<=0;
   22372: out<=0;
   22373: out<=1;
   22374: out<=0;
   22375: out<=1;
   22376: out<=0;
   22377: out<=1;
   22378: out<=1;
   22379: out<=0;
   22380: out<=1;
   22381: out<=1;
   22382: out<=1;
   22383: out<=1;
   22384: out<=1;
   22385: out<=1;
   22386: out<=0;
   22387: out<=0;
   22388: out<=0;
   22389: out<=1;
   22390: out<=0;
   22391: out<=1;
   22392: out<=0;
   22393: out<=1;
   22394: out<=1;
   22395: out<=0;
   22396: out<=1;
   22397: out<=1;
   22398: out<=1;
   22399: out<=1;
   22400: out<=0;
   22401: out<=0;
   22402: out<=1;
   22403: out<=1;
   22404: out<=1;
   22405: out<=0;
   22406: out<=1;
   22407: out<=0;
   22408: out<=1;
   22409: out<=0;
   22410: out<=0;
   22411: out<=1;
   22412: out<=0;
   22413: out<=0;
   22414: out<=0;
   22415: out<=0;
   22416: out<=0;
   22417: out<=0;
   22418: out<=1;
   22419: out<=1;
   22420: out<=1;
   22421: out<=0;
   22422: out<=1;
   22423: out<=0;
   22424: out<=1;
   22425: out<=0;
   22426: out<=0;
   22427: out<=1;
   22428: out<=0;
   22429: out<=0;
   22430: out<=0;
   22431: out<=0;
   22432: out<=1;
   22433: out<=1;
   22434: out<=0;
   22435: out<=0;
   22436: out<=0;
   22437: out<=1;
   22438: out<=0;
   22439: out<=1;
   22440: out<=0;
   22441: out<=1;
   22442: out<=1;
   22443: out<=0;
   22444: out<=1;
   22445: out<=1;
   22446: out<=1;
   22447: out<=1;
   22448: out<=1;
   22449: out<=1;
   22450: out<=0;
   22451: out<=0;
   22452: out<=0;
   22453: out<=1;
   22454: out<=0;
   22455: out<=1;
   22456: out<=0;
   22457: out<=1;
   22458: out<=1;
   22459: out<=0;
   22460: out<=1;
   22461: out<=1;
   22462: out<=1;
   22463: out<=1;
   22464: out<=0;
   22465: out<=0;
   22466: out<=1;
   22467: out<=1;
   22468: out<=1;
   22469: out<=0;
   22470: out<=1;
   22471: out<=0;
   22472: out<=1;
   22473: out<=0;
   22474: out<=0;
   22475: out<=1;
   22476: out<=0;
   22477: out<=0;
   22478: out<=0;
   22479: out<=0;
   22480: out<=1;
   22481: out<=1;
   22482: out<=0;
   22483: out<=0;
   22484: out<=0;
   22485: out<=1;
   22486: out<=0;
   22487: out<=1;
   22488: out<=0;
   22489: out<=1;
   22490: out<=1;
   22491: out<=0;
   22492: out<=1;
   22493: out<=1;
   22494: out<=1;
   22495: out<=1;
   22496: out<=0;
   22497: out<=0;
   22498: out<=1;
   22499: out<=1;
   22500: out<=1;
   22501: out<=0;
   22502: out<=1;
   22503: out<=0;
   22504: out<=1;
   22505: out<=0;
   22506: out<=0;
   22507: out<=1;
   22508: out<=0;
   22509: out<=0;
   22510: out<=0;
   22511: out<=0;
   22512: out<=1;
   22513: out<=1;
   22514: out<=0;
   22515: out<=0;
   22516: out<=0;
   22517: out<=1;
   22518: out<=0;
   22519: out<=1;
   22520: out<=0;
   22521: out<=1;
   22522: out<=1;
   22523: out<=0;
   22524: out<=1;
   22525: out<=1;
   22526: out<=1;
   22527: out<=1;
   22528: out<=1;
   22529: out<=1;
   22530: out<=0;
   22531: out<=0;
   22532: out<=0;
   22533: out<=1;
   22534: out<=0;
   22535: out<=1;
   22536: out<=1;
   22537: out<=0;
   22538: out<=0;
   22539: out<=1;
   22540: out<=0;
   22541: out<=0;
   22542: out<=0;
   22543: out<=0;
   22544: out<=0;
   22545: out<=0;
   22546: out<=1;
   22547: out<=1;
   22548: out<=1;
   22549: out<=0;
   22550: out<=1;
   22551: out<=0;
   22552: out<=0;
   22553: out<=1;
   22554: out<=1;
   22555: out<=0;
   22556: out<=1;
   22557: out<=1;
   22558: out<=1;
   22559: out<=1;
   22560: out<=1;
   22561: out<=1;
   22562: out<=0;
   22563: out<=0;
   22564: out<=0;
   22565: out<=1;
   22566: out<=0;
   22567: out<=1;
   22568: out<=1;
   22569: out<=0;
   22570: out<=0;
   22571: out<=1;
   22572: out<=0;
   22573: out<=0;
   22574: out<=0;
   22575: out<=0;
   22576: out<=0;
   22577: out<=0;
   22578: out<=1;
   22579: out<=1;
   22580: out<=1;
   22581: out<=0;
   22582: out<=1;
   22583: out<=0;
   22584: out<=0;
   22585: out<=1;
   22586: out<=1;
   22587: out<=0;
   22588: out<=1;
   22589: out<=1;
   22590: out<=1;
   22591: out<=1;
   22592: out<=1;
   22593: out<=1;
   22594: out<=0;
   22595: out<=0;
   22596: out<=0;
   22597: out<=1;
   22598: out<=0;
   22599: out<=1;
   22600: out<=1;
   22601: out<=0;
   22602: out<=0;
   22603: out<=1;
   22604: out<=0;
   22605: out<=0;
   22606: out<=0;
   22607: out<=0;
   22608: out<=1;
   22609: out<=1;
   22610: out<=0;
   22611: out<=0;
   22612: out<=0;
   22613: out<=1;
   22614: out<=0;
   22615: out<=1;
   22616: out<=1;
   22617: out<=0;
   22618: out<=0;
   22619: out<=1;
   22620: out<=0;
   22621: out<=0;
   22622: out<=0;
   22623: out<=0;
   22624: out<=0;
   22625: out<=0;
   22626: out<=1;
   22627: out<=1;
   22628: out<=1;
   22629: out<=0;
   22630: out<=1;
   22631: out<=0;
   22632: out<=0;
   22633: out<=1;
   22634: out<=1;
   22635: out<=0;
   22636: out<=1;
   22637: out<=1;
   22638: out<=1;
   22639: out<=1;
   22640: out<=0;
   22641: out<=0;
   22642: out<=1;
   22643: out<=1;
   22644: out<=1;
   22645: out<=0;
   22646: out<=1;
   22647: out<=0;
   22648: out<=0;
   22649: out<=1;
   22650: out<=1;
   22651: out<=0;
   22652: out<=1;
   22653: out<=1;
   22654: out<=1;
   22655: out<=1;
   22656: out<=0;
   22657: out<=0;
   22658: out<=1;
   22659: out<=1;
   22660: out<=1;
   22661: out<=0;
   22662: out<=1;
   22663: out<=0;
   22664: out<=0;
   22665: out<=1;
   22666: out<=1;
   22667: out<=0;
   22668: out<=1;
   22669: out<=1;
   22670: out<=1;
   22671: out<=1;
   22672: out<=0;
   22673: out<=0;
   22674: out<=1;
   22675: out<=1;
   22676: out<=1;
   22677: out<=0;
   22678: out<=1;
   22679: out<=0;
   22680: out<=0;
   22681: out<=1;
   22682: out<=1;
   22683: out<=0;
   22684: out<=1;
   22685: out<=1;
   22686: out<=1;
   22687: out<=1;
   22688: out<=0;
   22689: out<=0;
   22690: out<=1;
   22691: out<=1;
   22692: out<=1;
   22693: out<=0;
   22694: out<=1;
   22695: out<=0;
   22696: out<=0;
   22697: out<=1;
   22698: out<=1;
   22699: out<=0;
   22700: out<=1;
   22701: out<=1;
   22702: out<=1;
   22703: out<=1;
   22704: out<=0;
   22705: out<=0;
   22706: out<=1;
   22707: out<=1;
   22708: out<=1;
   22709: out<=0;
   22710: out<=1;
   22711: out<=0;
   22712: out<=0;
   22713: out<=1;
   22714: out<=1;
   22715: out<=0;
   22716: out<=1;
   22717: out<=1;
   22718: out<=1;
   22719: out<=1;
   22720: out<=0;
   22721: out<=0;
   22722: out<=1;
   22723: out<=1;
   22724: out<=1;
   22725: out<=0;
   22726: out<=1;
   22727: out<=0;
   22728: out<=0;
   22729: out<=1;
   22730: out<=1;
   22731: out<=0;
   22732: out<=1;
   22733: out<=1;
   22734: out<=1;
   22735: out<=1;
   22736: out<=1;
   22737: out<=1;
   22738: out<=0;
   22739: out<=0;
   22740: out<=0;
   22741: out<=1;
   22742: out<=0;
   22743: out<=1;
   22744: out<=1;
   22745: out<=0;
   22746: out<=0;
   22747: out<=1;
   22748: out<=0;
   22749: out<=0;
   22750: out<=0;
   22751: out<=0;
   22752: out<=1;
   22753: out<=1;
   22754: out<=0;
   22755: out<=0;
   22756: out<=0;
   22757: out<=1;
   22758: out<=0;
   22759: out<=1;
   22760: out<=1;
   22761: out<=0;
   22762: out<=0;
   22763: out<=1;
   22764: out<=0;
   22765: out<=0;
   22766: out<=0;
   22767: out<=0;
   22768: out<=0;
   22769: out<=0;
   22770: out<=1;
   22771: out<=1;
   22772: out<=1;
   22773: out<=0;
   22774: out<=1;
   22775: out<=0;
   22776: out<=0;
   22777: out<=1;
   22778: out<=1;
   22779: out<=0;
   22780: out<=1;
   22781: out<=1;
   22782: out<=1;
   22783: out<=1;
   22784: out<=0;
   22785: out<=1;
   22786: out<=0;
   22787: out<=1;
   22788: out<=0;
   22789: out<=0;
   22790: out<=1;
   22791: out<=1;
   22792: out<=1;
   22793: out<=1;
   22794: out<=1;
   22795: out<=1;
   22796: out<=1;
   22797: out<=0;
   22798: out<=0;
   22799: out<=1;
   22800: out<=0;
   22801: out<=1;
   22802: out<=0;
   22803: out<=1;
   22804: out<=0;
   22805: out<=0;
   22806: out<=1;
   22807: out<=1;
   22808: out<=1;
   22809: out<=1;
   22810: out<=1;
   22811: out<=1;
   22812: out<=1;
   22813: out<=0;
   22814: out<=0;
   22815: out<=1;
   22816: out<=1;
   22817: out<=0;
   22818: out<=1;
   22819: out<=0;
   22820: out<=1;
   22821: out<=1;
   22822: out<=0;
   22823: out<=0;
   22824: out<=0;
   22825: out<=0;
   22826: out<=0;
   22827: out<=0;
   22828: out<=0;
   22829: out<=1;
   22830: out<=1;
   22831: out<=0;
   22832: out<=1;
   22833: out<=0;
   22834: out<=1;
   22835: out<=0;
   22836: out<=1;
   22837: out<=1;
   22838: out<=0;
   22839: out<=0;
   22840: out<=0;
   22841: out<=0;
   22842: out<=0;
   22843: out<=0;
   22844: out<=0;
   22845: out<=1;
   22846: out<=1;
   22847: out<=0;
   22848: out<=0;
   22849: out<=1;
   22850: out<=0;
   22851: out<=1;
   22852: out<=0;
   22853: out<=0;
   22854: out<=1;
   22855: out<=1;
   22856: out<=1;
   22857: out<=1;
   22858: out<=1;
   22859: out<=1;
   22860: out<=1;
   22861: out<=0;
   22862: out<=0;
   22863: out<=1;
   22864: out<=1;
   22865: out<=0;
   22866: out<=1;
   22867: out<=0;
   22868: out<=1;
   22869: out<=1;
   22870: out<=0;
   22871: out<=0;
   22872: out<=0;
   22873: out<=0;
   22874: out<=0;
   22875: out<=0;
   22876: out<=0;
   22877: out<=1;
   22878: out<=1;
   22879: out<=0;
   22880: out<=0;
   22881: out<=1;
   22882: out<=0;
   22883: out<=1;
   22884: out<=0;
   22885: out<=0;
   22886: out<=1;
   22887: out<=1;
   22888: out<=1;
   22889: out<=1;
   22890: out<=1;
   22891: out<=1;
   22892: out<=1;
   22893: out<=0;
   22894: out<=0;
   22895: out<=1;
   22896: out<=1;
   22897: out<=0;
   22898: out<=1;
   22899: out<=0;
   22900: out<=1;
   22901: out<=1;
   22902: out<=0;
   22903: out<=0;
   22904: out<=0;
   22905: out<=0;
   22906: out<=0;
   22907: out<=0;
   22908: out<=0;
   22909: out<=1;
   22910: out<=1;
   22911: out<=0;
   22912: out<=1;
   22913: out<=0;
   22914: out<=1;
   22915: out<=0;
   22916: out<=1;
   22917: out<=1;
   22918: out<=0;
   22919: out<=0;
   22920: out<=0;
   22921: out<=0;
   22922: out<=0;
   22923: out<=0;
   22924: out<=0;
   22925: out<=1;
   22926: out<=1;
   22927: out<=0;
   22928: out<=0;
   22929: out<=1;
   22930: out<=0;
   22931: out<=1;
   22932: out<=0;
   22933: out<=0;
   22934: out<=1;
   22935: out<=1;
   22936: out<=1;
   22937: out<=1;
   22938: out<=1;
   22939: out<=1;
   22940: out<=1;
   22941: out<=0;
   22942: out<=0;
   22943: out<=1;
   22944: out<=0;
   22945: out<=1;
   22946: out<=0;
   22947: out<=1;
   22948: out<=0;
   22949: out<=0;
   22950: out<=1;
   22951: out<=1;
   22952: out<=1;
   22953: out<=1;
   22954: out<=1;
   22955: out<=1;
   22956: out<=1;
   22957: out<=0;
   22958: out<=0;
   22959: out<=1;
   22960: out<=1;
   22961: out<=0;
   22962: out<=1;
   22963: out<=0;
   22964: out<=1;
   22965: out<=1;
   22966: out<=0;
   22967: out<=0;
   22968: out<=0;
   22969: out<=0;
   22970: out<=0;
   22971: out<=0;
   22972: out<=0;
   22973: out<=1;
   22974: out<=1;
   22975: out<=0;
   22976: out<=1;
   22977: out<=0;
   22978: out<=1;
   22979: out<=0;
   22980: out<=1;
   22981: out<=1;
   22982: out<=0;
   22983: out<=0;
   22984: out<=0;
   22985: out<=0;
   22986: out<=0;
   22987: out<=0;
   22988: out<=0;
   22989: out<=1;
   22990: out<=1;
   22991: out<=0;
   22992: out<=1;
   22993: out<=0;
   22994: out<=1;
   22995: out<=0;
   22996: out<=1;
   22997: out<=1;
   22998: out<=0;
   22999: out<=0;
   23000: out<=0;
   23001: out<=0;
   23002: out<=0;
   23003: out<=0;
   23004: out<=0;
   23005: out<=1;
   23006: out<=1;
   23007: out<=0;
   23008: out<=1;
   23009: out<=0;
   23010: out<=1;
   23011: out<=0;
   23012: out<=1;
   23013: out<=1;
   23014: out<=0;
   23015: out<=0;
   23016: out<=0;
   23017: out<=0;
   23018: out<=0;
   23019: out<=0;
   23020: out<=0;
   23021: out<=1;
   23022: out<=1;
   23023: out<=0;
   23024: out<=1;
   23025: out<=0;
   23026: out<=1;
   23027: out<=0;
   23028: out<=1;
   23029: out<=1;
   23030: out<=0;
   23031: out<=0;
   23032: out<=0;
   23033: out<=0;
   23034: out<=0;
   23035: out<=0;
   23036: out<=0;
   23037: out<=1;
   23038: out<=1;
   23039: out<=0;
   23040: out<=1;
   23041: out<=0;
   23042: out<=0;
   23043: out<=1;
   23044: out<=1;
   23045: out<=1;
   23046: out<=1;
   23047: out<=1;
   23048: out<=1;
   23049: out<=1;
   23050: out<=0;
   23051: out<=0;
   23052: out<=1;
   23053: out<=0;
   23054: out<=1;
   23055: out<=0;
   23056: out<=1;
   23057: out<=0;
   23058: out<=0;
   23059: out<=1;
   23060: out<=1;
   23061: out<=1;
   23062: out<=1;
   23063: out<=1;
   23064: out<=1;
   23065: out<=1;
   23066: out<=0;
   23067: out<=0;
   23068: out<=1;
   23069: out<=0;
   23070: out<=1;
   23071: out<=0;
   23072: out<=1;
   23073: out<=0;
   23074: out<=0;
   23075: out<=1;
   23076: out<=1;
   23077: out<=1;
   23078: out<=1;
   23079: out<=1;
   23080: out<=1;
   23081: out<=1;
   23082: out<=0;
   23083: out<=0;
   23084: out<=1;
   23085: out<=0;
   23086: out<=1;
   23087: out<=0;
   23088: out<=1;
   23089: out<=0;
   23090: out<=0;
   23091: out<=1;
   23092: out<=1;
   23093: out<=1;
   23094: out<=1;
   23095: out<=1;
   23096: out<=1;
   23097: out<=1;
   23098: out<=0;
   23099: out<=0;
   23100: out<=1;
   23101: out<=0;
   23102: out<=1;
   23103: out<=0;
   23104: out<=1;
   23105: out<=0;
   23106: out<=0;
   23107: out<=1;
   23108: out<=1;
   23109: out<=1;
   23110: out<=1;
   23111: out<=1;
   23112: out<=1;
   23113: out<=1;
   23114: out<=0;
   23115: out<=0;
   23116: out<=1;
   23117: out<=0;
   23118: out<=1;
   23119: out<=0;
   23120: out<=0;
   23121: out<=1;
   23122: out<=1;
   23123: out<=0;
   23124: out<=0;
   23125: out<=0;
   23126: out<=0;
   23127: out<=0;
   23128: out<=0;
   23129: out<=0;
   23130: out<=1;
   23131: out<=1;
   23132: out<=0;
   23133: out<=1;
   23134: out<=0;
   23135: out<=1;
   23136: out<=0;
   23137: out<=1;
   23138: out<=1;
   23139: out<=0;
   23140: out<=0;
   23141: out<=0;
   23142: out<=0;
   23143: out<=0;
   23144: out<=0;
   23145: out<=0;
   23146: out<=1;
   23147: out<=1;
   23148: out<=0;
   23149: out<=1;
   23150: out<=0;
   23151: out<=1;
   23152: out<=1;
   23153: out<=0;
   23154: out<=0;
   23155: out<=1;
   23156: out<=1;
   23157: out<=1;
   23158: out<=1;
   23159: out<=1;
   23160: out<=1;
   23161: out<=1;
   23162: out<=0;
   23163: out<=0;
   23164: out<=1;
   23165: out<=0;
   23166: out<=1;
   23167: out<=0;
   23168: out<=0;
   23169: out<=1;
   23170: out<=1;
   23171: out<=0;
   23172: out<=0;
   23173: out<=0;
   23174: out<=0;
   23175: out<=0;
   23176: out<=0;
   23177: out<=0;
   23178: out<=1;
   23179: out<=1;
   23180: out<=0;
   23181: out<=1;
   23182: out<=0;
   23183: out<=1;
   23184: out<=1;
   23185: out<=0;
   23186: out<=0;
   23187: out<=1;
   23188: out<=1;
   23189: out<=1;
   23190: out<=1;
   23191: out<=1;
   23192: out<=1;
   23193: out<=1;
   23194: out<=0;
   23195: out<=0;
   23196: out<=1;
   23197: out<=0;
   23198: out<=1;
   23199: out<=0;
   23200: out<=0;
   23201: out<=1;
   23202: out<=1;
   23203: out<=0;
   23204: out<=0;
   23205: out<=0;
   23206: out<=0;
   23207: out<=0;
   23208: out<=0;
   23209: out<=0;
   23210: out<=1;
   23211: out<=1;
   23212: out<=0;
   23213: out<=1;
   23214: out<=0;
   23215: out<=1;
   23216: out<=1;
   23217: out<=0;
   23218: out<=0;
   23219: out<=1;
   23220: out<=1;
   23221: out<=1;
   23222: out<=1;
   23223: out<=1;
   23224: out<=1;
   23225: out<=1;
   23226: out<=0;
   23227: out<=0;
   23228: out<=1;
   23229: out<=0;
   23230: out<=1;
   23231: out<=0;
   23232: out<=0;
   23233: out<=1;
   23234: out<=1;
   23235: out<=0;
   23236: out<=0;
   23237: out<=0;
   23238: out<=0;
   23239: out<=0;
   23240: out<=0;
   23241: out<=0;
   23242: out<=1;
   23243: out<=1;
   23244: out<=0;
   23245: out<=1;
   23246: out<=0;
   23247: out<=1;
   23248: out<=0;
   23249: out<=1;
   23250: out<=1;
   23251: out<=0;
   23252: out<=0;
   23253: out<=0;
   23254: out<=0;
   23255: out<=0;
   23256: out<=0;
   23257: out<=0;
   23258: out<=1;
   23259: out<=1;
   23260: out<=0;
   23261: out<=1;
   23262: out<=0;
   23263: out<=1;
   23264: out<=1;
   23265: out<=0;
   23266: out<=0;
   23267: out<=1;
   23268: out<=1;
   23269: out<=1;
   23270: out<=1;
   23271: out<=1;
   23272: out<=1;
   23273: out<=1;
   23274: out<=0;
   23275: out<=0;
   23276: out<=1;
   23277: out<=0;
   23278: out<=1;
   23279: out<=0;
   23280: out<=1;
   23281: out<=0;
   23282: out<=0;
   23283: out<=1;
   23284: out<=1;
   23285: out<=1;
   23286: out<=1;
   23287: out<=1;
   23288: out<=1;
   23289: out<=1;
   23290: out<=0;
   23291: out<=0;
   23292: out<=1;
   23293: out<=0;
   23294: out<=1;
   23295: out<=0;
   23296: out<=0;
   23297: out<=0;
   23298: out<=0;
   23299: out<=0;
   23300: out<=1;
   23301: out<=0;
   23302: out<=0;
   23303: out<=1;
   23304: out<=1;
   23305: out<=0;
   23306: out<=1;
   23307: out<=0;
   23308: out<=0;
   23309: out<=0;
   23310: out<=1;
   23311: out<=1;
   23312: out<=1;
   23313: out<=1;
   23314: out<=1;
   23315: out<=1;
   23316: out<=0;
   23317: out<=1;
   23318: out<=1;
   23319: out<=0;
   23320: out<=0;
   23321: out<=1;
   23322: out<=0;
   23323: out<=1;
   23324: out<=1;
   23325: out<=1;
   23326: out<=0;
   23327: out<=0;
   23328: out<=1;
   23329: out<=1;
   23330: out<=1;
   23331: out<=1;
   23332: out<=0;
   23333: out<=1;
   23334: out<=1;
   23335: out<=0;
   23336: out<=0;
   23337: out<=1;
   23338: out<=0;
   23339: out<=1;
   23340: out<=1;
   23341: out<=1;
   23342: out<=0;
   23343: out<=0;
   23344: out<=0;
   23345: out<=0;
   23346: out<=0;
   23347: out<=0;
   23348: out<=1;
   23349: out<=0;
   23350: out<=0;
   23351: out<=1;
   23352: out<=1;
   23353: out<=0;
   23354: out<=1;
   23355: out<=0;
   23356: out<=0;
   23357: out<=0;
   23358: out<=1;
   23359: out<=1;
   23360: out<=0;
   23361: out<=0;
   23362: out<=0;
   23363: out<=0;
   23364: out<=1;
   23365: out<=0;
   23366: out<=0;
   23367: out<=1;
   23368: out<=1;
   23369: out<=0;
   23370: out<=1;
   23371: out<=0;
   23372: out<=0;
   23373: out<=0;
   23374: out<=1;
   23375: out<=1;
   23376: out<=0;
   23377: out<=0;
   23378: out<=0;
   23379: out<=0;
   23380: out<=1;
   23381: out<=0;
   23382: out<=0;
   23383: out<=1;
   23384: out<=1;
   23385: out<=0;
   23386: out<=1;
   23387: out<=0;
   23388: out<=0;
   23389: out<=0;
   23390: out<=1;
   23391: out<=1;
   23392: out<=0;
   23393: out<=0;
   23394: out<=0;
   23395: out<=0;
   23396: out<=1;
   23397: out<=0;
   23398: out<=0;
   23399: out<=1;
   23400: out<=1;
   23401: out<=0;
   23402: out<=1;
   23403: out<=0;
   23404: out<=0;
   23405: out<=0;
   23406: out<=1;
   23407: out<=1;
   23408: out<=0;
   23409: out<=0;
   23410: out<=0;
   23411: out<=0;
   23412: out<=1;
   23413: out<=0;
   23414: out<=0;
   23415: out<=1;
   23416: out<=1;
   23417: out<=0;
   23418: out<=1;
   23419: out<=0;
   23420: out<=0;
   23421: out<=0;
   23422: out<=1;
   23423: out<=1;
   23424: out<=1;
   23425: out<=1;
   23426: out<=1;
   23427: out<=1;
   23428: out<=0;
   23429: out<=1;
   23430: out<=1;
   23431: out<=0;
   23432: out<=0;
   23433: out<=1;
   23434: out<=0;
   23435: out<=1;
   23436: out<=1;
   23437: out<=1;
   23438: out<=0;
   23439: out<=0;
   23440: out<=1;
   23441: out<=1;
   23442: out<=1;
   23443: out<=1;
   23444: out<=0;
   23445: out<=1;
   23446: out<=1;
   23447: out<=0;
   23448: out<=0;
   23449: out<=1;
   23450: out<=0;
   23451: out<=1;
   23452: out<=1;
   23453: out<=1;
   23454: out<=0;
   23455: out<=0;
   23456: out<=0;
   23457: out<=0;
   23458: out<=0;
   23459: out<=0;
   23460: out<=1;
   23461: out<=0;
   23462: out<=0;
   23463: out<=1;
   23464: out<=1;
   23465: out<=0;
   23466: out<=1;
   23467: out<=0;
   23468: out<=0;
   23469: out<=0;
   23470: out<=1;
   23471: out<=1;
   23472: out<=0;
   23473: out<=0;
   23474: out<=0;
   23475: out<=0;
   23476: out<=1;
   23477: out<=0;
   23478: out<=0;
   23479: out<=1;
   23480: out<=1;
   23481: out<=0;
   23482: out<=1;
   23483: out<=0;
   23484: out<=0;
   23485: out<=0;
   23486: out<=1;
   23487: out<=1;
   23488: out<=1;
   23489: out<=1;
   23490: out<=1;
   23491: out<=1;
   23492: out<=0;
   23493: out<=1;
   23494: out<=1;
   23495: out<=0;
   23496: out<=0;
   23497: out<=1;
   23498: out<=0;
   23499: out<=1;
   23500: out<=1;
   23501: out<=1;
   23502: out<=0;
   23503: out<=0;
   23504: out<=0;
   23505: out<=0;
   23506: out<=0;
   23507: out<=0;
   23508: out<=1;
   23509: out<=0;
   23510: out<=0;
   23511: out<=1;
   23512: out<=1;
   23513: out<=0;
   23514: out<=1;
   23515: out<=0;
   23516: out<=0;
   23517: out<=0;
   23518: out<=1;
   23519: out<=1;
   23520: out<=1;
   23521: out<=1;
   23522: out<=1;
   23523: out<=1;
   23524: out<=0;
   23525: out<=1;
   23526: out<=1;
   23527: out<=0;
   23528: out<=0;
   23529: out<=1;
   23530: out<=0;
   23531: out<=1;
   23532: out<=1;
   23533: out<=1;
   23534: out<=0;
   23535: out<=0;
   23536: out<=0;
   23537: out<=0;
   23538: out<=0;
   23539: out<=0;
   23540: out<=1;
   23541: out<=0;
   23542: out<=0;
   23543: out<=1;
   23544: out<=1;
   23545: out<=0;
   23546: out<=1;
   23547: out<=0;
   23548: out<=0;
   23549: out<=0;
   23550: out<=1;
   23551: out<=1;
   23552: out<=1;
   23553: out<=0;
   23554: out<=1;
   23555: out<=0;
   23556: out<=0;
   23557: out<=0;
   23558: out<=1;
   23559: out<=1;
   23560: out<=1;
   23561: out<=1;
   23562: out<=1;
   23563: out<=1;
   23564: out<=0;
   23565: out<=1;
   23566: out<=1;
   23567: out<=0;
   23568: out<=0;
   23569: out<=1;
   23570: out<=0;
   23571: out<=1;
   23572: out<=1;
   23573: out<=1;
   23574: out<=0;
   23575: out<=0;
   23576: out<=0;
   23577: out<=0;
   23578: out<=0;
   23579: out<=0;
   23580: out<=1;
   23581: out<=0;
   23582: out<=0;
   23583: out<=1;
   23584: out<=1;
   23585: out<=0;
   23586: out<=1;
   23587: out<=0;
   23588: out<=0;
   23589: out<=0;
   23590: out<=1;
   23591: out<=1;
   23592: out<=1;
   23593: out<=1;
   23594: out<=1;
   23595: out<=1;
   23596: out<=0;
   23597: out<=1;
   23598: out<=1;
   23599: out<=0;
   23600: out<=0;
   23601: out<=1;
   23602: out<=0;
   23603: out<=1;
   23604: out<=1;
   23605: out<=1;
   23606: out<=0;
   23607: out<=0;
   23608: out<=0;
   23609: out<=0;
   23610: out<=0;
   23611: out<=0;
   23612: out<=1;
   23613: out<=0;
   23614: out<=0;
   23615: out<=1;
   23616: out<=1;
   23617: out<=0;
   23618: out<=1;
   23619: out<=0;
   23620: out<=0;
   23621: out<=0;
   23622: out<=1;
   23623: out<=1;
   23624: out<=1;
   23625: out<=1;
   23626: out<=1;
   23627: out<=1;
   23628: out<=0;
   23629: out<=1;
   23630: out<=1;
   23631: out<=0;
   23632: out<=1;
   23633: out<=0;
   23634: out<=1;
   23635: out<=0;
   23636: out<=0;
   23637: out<=0;
   23638: out<=1;
   23639: out<=1;
   23640: out<=1;
   23641: out<=1;
   23642: out<=1;
   23643: out<=1;
   23644: out<=0;
   23645: out<=1;
   23646: out<=1;
   23647: out<=0;
   23648: out<=0;
   23649: out<=1;
   23650: out<=0;
   23651: out<=1;
   23652: out<=1;
   23653: out<=1;
   23654: out<=0;
   23655: out<=0;
   23656: out<=0;
   23657: out<=0;
   23658: out<=0;
   23659: out<=0;
   23660: out<=1;
   23661: out<=0;
   23662: out<=0;
   23663: out<=1;
   23664: out<=0;
   23665: out<=1;
   23666: out<=0;
   23667: out<=1;
   23668: out<=1;
   23669: out<=1;
   23670: out<=0;
   23671: out<=0;
   23672: out<=0;
   23673: out<=0;
   23674: out<=0;
   23675: out<=0;
   23676: out<=1;
   23677: out<=0;
   23678: out<=0;
   23679: out<=1;
   23680: out<=0;
   23681: out<=1;
   23682: out<=0;
   23683: out<=1;
   23684: out<=1;
   23685: out<=1;
   23686: out<=0;
   23687: out<=0;
   23688: out<=0;
   23689: out<=0;
   23690: out<=0;
   23691: out<=0;
   23692: out<=1;
   23693: out<=0;
   23694: out<=0;
   23695: out<=1;
   23696: out<=0;
   23697: out<=1;
   23698: out<=0;
   23699: out<=1;
   23700: out<=1;
   23701: out<=1;
   23702: out<=0;
   23703: out<=0;
   23704: out<=0;
   23705: out<=0;
   23706: out<=0;
   23707: out<=0;
   23708: out<=1;
   23709: out<=0;
   23710: out<=0;
   23711: out<=1;
   23712: out<=0;
   23713: out<=1;
   23714: out<=0;
   23715: out<=1;
   23716: out<=1;
   23717: out<=1;
   23718: out<=0;
   23719: out<=0;
   23720: out<=0;
   23721: out<=0;
   23722: out<=0;
   23723: out<=0;
   23724: out<=1;
   23725: out<=0;
   23726: out<=0;
   23727: out<=1;
   23728: out<=0;
   23729: out<=1;
   23730: out<=0;
   23731: out<=1;
   23732: out<=1;
   23733: out<=1;
   23734: out<=0;
   23735: out<=0;
   23736: out<=0;
   23737: out<=0;
   23738: out<=0;
   23739: out<=0;
   23740: out<=1;
   23741: out<=0;
   23742: out<=0;
   23743: out<=1;
   23744: out<=0;
   23745: out<=1;
   23746: out<=0;
   23747: out<=1;
   23748: out<=1;
   23749: out<=1;
   23750: out<=0;
   23751: out<=0;
   23752: out<=0;
   23753: out<=0;
   23754: out<=0;
   23755: out<=0;
   23756: out<=1;
   23757: out<=0;
   23758: out<=0;
   23759: out<=1;
   23760: out<=1;
   23761: out<=0;
   23762: out<=1;
   23763: out<=0;
   23764: out<=0;
   23765: out<=0;
   23766: out<=1;
   23767: out<=1;
   23768: out<=1;
   23769: out<=1;
   23770: out<=1;
   23771: out<=1;
   23772: out<=0;
   23773: out<=1;
   23774: out<=1;
   23775: out<=0;
   23776: out<=1;
   23777: out<=0;
   23778: out<=1;
   23779: out<=0;
   23780: out<=0;
   23781: out<=0;
   23782: out<=1;
   23783: out<=1;
   23784: out<=1;
   23785: out<=1;
   23786: out<=1;
   23787: out<=1;
   23788: out<=0;
   23789: out<=1;
   23790: out<=1;
   23791: out<=0;
   23792: out<=0;
   23793: out<=1;
   23794: out<=0;
   23795: out<=1;
   23796: out<=1;
   23797: out<=1;
   23798: out<=0;
   23799: out<=0;
   23800: out<=0;
   23801: out<=0;
   23802: out<=0;
   23803: out<=0;
   23804: out<=1;
   23805: out<=0;
   23806: out<=0;
   23807: out<=1;
   23808: out<=1;
   23809: out<=1;
   23810: out<=0;
   23811: out<=0;
   23812: out<=1;
   23813: out<=0;
   23814: out<=1;
   23815: out<=0;
   23816: out<=0;
   23817: out<=1;
   23818: out<=1;
   23819: out<=0;
   23820: out<=0;
   23821: out<=0;
   23822: out<=0;
   23823: out<=0;
   23824: out<=1;
   23825: out<=1;
   23826: out<=0;
   23827: out<=0;
   23828: out<=1;
   23829: out<=0;
   23830: out<=1;
   23831: out<=0;
   23832: out<=0;
   23833: out<=1;
   23834: out<=1;
   23835: out<=0;
   23836: out<=0;
   23837: out<=0;
   23838: out<=0;
   23839: out<=0;
   23840: out<=0;
   23841: out<=0;
   23842: out<=1;
   23843: out<=1;
   23844: out<=0;
   23845: out<=1;
   23846: out<=0;
   23847: out<=1;
   23848: out<=1;
   23849: out<=0;
   23850: out<=0;
   23851: out<=1;
   23852: out<=1;
   23853: out<=1;
   23854: out<=1;
   23855: out<=1;
   23856: out<=0;
   23857: out<=0;
   23858: out<=1;
   23859: out<=1;
   23860: out<=0;
   23861: out<=1;
   23862: out<=0;
   23863: out<=1;
   23864: out<=1;
   23865: out<=0;
   23866: out<=0;
   23867: out<=1;
   23868: out<=1;
   23869: out<=1;
   23870: out<=1;
   23871: out<=1;
   23872: out<=1;
   23873: out<=1;
   23874: out<=0;
   23875: out<=0;
   23876: out<=1;
   23877: out<=0;
   23878: out<=1;
   23879: out<=0;
   23880: out<=0;
   23881: out<=1;
   23882: out<=1;
   23883: out<=0;
   23884: out<=0;
   23885: out<=0;
   23886: out<=0;
   23887: out<=0;
   23888: out<=0;
   23889: out<=0;
   23890: out<=1;
   23891: out<=1;
   23892: out<=0;
   23893: out<=1;
   23894: out<=0;
   23895: out<=1;
   23896: out<=1;
   23897: out<=0;
   23898: out<=0;
   23899: out<=1;
   23900: out<=1;
   23901: out<=1;
   23902: out<=1;
   23903: out<=1;
   23904: out<=1;
   23905: out<=1;
   23906: out<=0;
   23907: out<=0;
   23908: out<=1;
   23909: out<=0;
   23910: out<=1;
   23911: out<=0;
   23912: out<=0;
   23913: out<=1;
   23914: out<=1;
   23915: out<=0;
   23916: out<=0;
   23917: out<=0;
   23918: out<=0;
   23919: out<=0;
   23920: out<=0;
   23921: out<=0;
   23922: out<=1;
   23923: out<=1;
   23924: out<=0;
   23925: out<=1;
   23926: out<=0;
   23927: out<=1;
   23928: out<=1;
   23929: out<=0;
   23930: out<=0;
   23931: out<=1;
   23932: out<=1;
   23933: out<=1;
   23934: out<=1;
   23935: out<=1;
   23936: out<=0;
   23937: out<=0;
   23938: out<=1;
   23939: out<=1;
   23940: out<=0;
   23941: out<=1;
   23942: out<=0;
   23943: out<=1;
   23944: out<=1;
   23945: out<=0;
   23946: out<=0;
   23947: out<=1;
   23948: out<=1;
   23949: out<=1;
   23950: out<=1;
   23951: out<=1;
   23952: out<=1;
   23953: out<=1;
   23954: out<=0;
   23955: out<=0;
   23956: out<=1;
   23957: out<=0;
   23958: out<=1;
   23959: out<=0;
   23960: out<=0;
   23961: out<=1;
   23962: out<=1;
   23963: out<=0;
   23964: out<=0;
   23965: out<=0;
   23966: out<=0;
   23967: out<=0;
   23968: out<=1;
   23969: out<=1;
   23970: out<=0;
   23971: out<=0;
   23972: out<=1;
   23973: out<=0;
   23974: out<=1;
   23975: out<=0;
   23976: out<=0;
   23977: out<=1;
   23978: out<=1;
   23979: out<=0;
   23980: out<=0;
   23981: out<=0;
   23982: out<=0;
   23983: out<=0;
   23984: out<=0;
   23985: out<=0;
   23986: out<=1;
   23987: out<=1;
   23988: out<=0;
   23989: out<=1;
   23990: out<=0;
   23991: out<=1;
   23992: out<=1;
   23993: out<=0;
   23994: out<=0;
   23995: out<=1;
   23996: out<=1;
   23997: out<=1;
   23998: out<=1;
   23999: out<=1;
   24000: out<=0;
   24001: out<=0;
   24002: out<=1;
   24003: out<=1;
   24004: out<=0;
   24005: out<=1;
   24006: out<=0;
   24007: out<=1;
   24008: out<=1;
   24009: out<=0;
   24010: out<=0;
   24011: out<=1;
   24012: out<=1;
   24013: out<=1;
   24014: out<=1;
   24015: out<=1;
   24016: out<=0;
   24017: out<=0;
   24018: out<=1;
   24019: out<=1;
   24020: out<=0;
   24021: out<=1;
   24022: out<=0;
   24023: out<=1;
   24024: out<=1;
   24025: out<=0;
   24026: out<=0;
   24027: out<=1;
   24028: out<=1;
   24029: out<=1;
   24030: out<=1;
   24031: out<=1;
   24032: out<=0;
   24033: out<=0;
   24034: out<=1;
   24035: out<=1;
   24036: out<=0;
   24037: out<=1;
   24038: out<=0;
   24039: out<=1;
   24040: out<=1;
   24041: out<=0;
   24042: out<=0;
   24043: out<=1;
   24044: out<=1;
   24045: out<=1;
   24046: out<=1;
   24047: out<=1;
   24048: out<=0;
   24049: out<=0;
   24050: out<=1;
   24051: out<=1;
   24052: out<=0;
   24053: out<=1;
   24054: out<=0;
   24055: out<=1;
   24056: out<=1;
   24057: out<=0;
   24058: out<=0;
   24059: out<=1;
   24060: out<=1;
   24061: out<=1;
   24062: out<=1;
   24063: out<=1;
   24064: out<=0;
   24065: out<=0;
   24066: out<=0;
   24067: out<=0;
   24068: out<=0;
   24069: out<=1;
   24070: out<=1;
   24071: out<=0;
   24072: out<=0;
   24073: out<=1;
   24074: out<=0;
   24075: out<=1;
   24076: out<=0;
   24077: out<=0;
   24078: out<=1;
   24079: out<=1;
   24080: out<=0;
   24081: out<=0;
   24082: out<=0;
   24083: out<=0;
   24084: out<=0;
   24085: out<=1;
   24086: out<=1;
   24087: out<=0;
   24088: out<=0;
   24089: out<=1;
   24090: out<=0;
   24091: out<=1;
   24092: out<=0;
   24093: out<=0;
   24094: out<=1;
   24095: out<=1;
   24096: out<=0;
   24097: out<=0;
   24098: out<=0;
   24099: out<=0;
   24100: out<=0;
   24101: out<=1;
   24102: out<=1;
   24103: out<=0;
   24104: out<=0;
   24105: out<=1;
   24106: out<=0;
   24107: out<=1;
   24108: out<=0;
   24109: out<=0;
   24110: out<=1;
   24111: out<=1;
   24112: out<=0;
   24113: out<=0;
   24114: out<=0;
   24115: out<=0;
   24116: out<=0;
   24117: out<=1;
   24118: out<=1;
   24119: out<=0;
   24120: out<=0;
   24121: out<=1;
   24122: out<=0;
   24123: out<=1;
   24124: out<=0;
   24125: out<=0;
   24126: out<=1;
   24127: out<=1;
   24128: out<=0;
   24129: out<=0;
   24130: out<=0;
   24131: out<=0;
   24132: out<=0;
   24133: out<=1;
   24134: out<=1;
   24135: out<=0;
   24136: out<=0;
   24137: out<=1;
   24138: out<=0;
   24139: out<=1;
   24140: out<=0;
   24141: out<=0;
   24142: out<=1;
   24143: out<=1;
   24144: out<=1;
   24145: out<=1;
   24146: out<=1;
   24147: out<=1;
   24148: out<=1;
   24149: out<=0;
   24150: out<=0;
   24151: out<=1;
   24152: out<=1;
   24153: out<=0;
   24154: out<=1;
   24155: out<=0;
   24156: out<=1;
   24157: out<=1;
   24158: out<=0;
   24159: out<=0;
   24160: out<=1;
   24161: out<=1;
   24162: out<=1;
   24163: out<=1;
   24164: out<=1;
   24165: out<=0;
   24166: out<=0;
   24167: out<=1;
   24168: out<=1;
   24169: out<=0;
   24170: out<=1;
   24171: out<=0;
   24172: out<=1;
   24173: out<=1;
   24174: out<=0;
   24175: out<=0;
   24176: out<=0;
   24177: out<=0;
   24178: out<=0;
   24179: out<=0;
   24180: out<=0;
   24181: out<=1;
   24182: out<=1;
   24183: out<=0;
   24184: out<=0;
   24185: out<=1;
   24186: out<=0;
   24187: out<=1;
   24188: out<=0;
   24189: out<=0;
   24190: out<=1;
   24191: out<=1;
   24192: out<=1;
   24193: out<=1;
   24194: out<=1;
   24195: out<=1;
   24196: out<=1;
   24197: out<=0;
   24198: out<=0;
   24199: out<=1;
   24200: out<=1;
   24201: out<=0;
   24202: out<=1;
   24203: out<=0;
   24204: out<=1;
   24205: out<=1;
   24206: out<=0;
   24207: out<=0;
   24208: out<=0;
   24209: out<=0;
   24210: out<=0;
   24211: out<=0;
   24212: out<=0;
   24213: out<=1;
   24214: out<=1;
   24215: out<=0;
   24216: out<=0;
   24217: out<=1;
   24218: out<=0;
   24219: out<=1;
   24220: out<=0;
   24221: out<=0;
   24222: out<=1;
   24223: out<=1;
   24224: out<=1;
   24225: out<=1;
   24226: out<=1;
   24227: out<=1;
   24228: out<=1;
   24229: out<=0;
   24230: out<=0;
   24231: out<=1;
   24232: out<=1;
   24233: out<=0;
   24234: out<=1;
   24235: out<=0;
   24236: out<=1;
   24237: out<=1;
   24238: out<=0;
   24239: out<=0;
   24240: out<=0;
   24241: out<=0;
   24242: out<=0;
   24243: out<=0;
   24244: out<=0;
   24245: out<=1;
   24246: out<=1;
   24247: out<=0;
   24248: out<=0;
   24249: out<=1;
   24250: out<=0;
   24251: out<=1;
   24252: out<=0;
   24253: out<=0;
   24254: out<=1;
   24255: out<=1;
   24256: out<=1;
   24257: out<=1;
   24258: out<=1;
   24259: out<=1;
   24260: out<=1;
   24261: out<=0;
   24262: out<=0;
   24263: out<=1;
   24264: out<=1;
   24265: out<=0;
   24266: out<=1;
   24267: out<=0;
   24268: out<=1;
   24269: out<=1;
   24270: out<=0;
   24271: out<=0;
   24272: out<=1;
   24273: out<=1;
   24274: out<=1;
   24275: out<=1;
   24276: out<=1;
   24277: out<=0;
   24278: out<=0;
   24279: out<=1;
   24280: out<=1;
   24281: out<=0;
   24282: out<=1;
   24283: out<=0;
   24284: out<=1;
   24285: out<=1;
   24286: out<=0;
   24287: out<=0;
   24288: out<=0;
   24289: out<=0;
   24290: out<=0;
   24291: out<=0;
   24292: out<=0;
   24293: out<=1;
   24294: out<=1;
   24295: out<=0;
   24296: out<=0;
   24297: out<=1;
   24298: out<=0;
   24299: out<=1;
   24300: out<=0;
   24301: out<=0;
   24302: out<=1;
   24303: out<=1;
   24304: out<=0;
   24305: out<=0;
   24306: out<=0;
   24307: out<=0;
   24308: out<=0;
   24309: out<=1;
   24310: out<=1;
   24311: out<=0;
   24312: out<=0;
   24313: out<=1;
   24314: out<=0;
   24315: out<=1;
   24316: out<=0;
   24317: out<=0;
   24318: out<=1;
   24319: out<=1;
   24320: out<=0;
   24321: out<=1;
   24322: out<=1;
   24323: out<=0;
   24324: out<=1;
   24325: out<=1;
   24326: out<=1;
   24327: out<=1;
   24328: out<=1;
   24329: out<=1;
   24330: out<=0;
   24331: out<=0;
   24332: out<=0;
   24333: out<=1;
   24334: out<=0;
   24335: out<=1;
   24336: out<=1;
   24337: out<=0;
   24338: out<=0;
   24339: out<=1;
   24340: out<=0;
   24341: out<=0;
   24342: out<=0;
   24343: out<=0;
   24344: out<=0;
   24345: out<=0;
   24346: out<=1;
   24347: out<=1;
   24348: out<=1;
   24349: out<=0;
   24350: out<=1;
   24351: out<=0;
   24352: out<=1;
   24353: out<=0;
   24354: out<=0;
   24355: out<=1;
   24356: out<=0;
   24357: out<=0;
   24358: out<=0;
   24359: out<=0;
   24360: out<=0;
   24361: out<=0;
   24362: out<=1;
   24363: out<=1;
   24364: out<=1;
   24365: out<=0;
   24366: out<=1;
   24367: out<=0;
   24368: out<=0;
   24369: out<=1;
   24370: out<=1;
   24371: out<=0;
   24372: out<=1;
   24373: out<=1;
   24374: out<=1;
   24375: out<=1;
   24376: out<=1;
   24377: out<=1;
   24378: out<=0;
   24379: out<=0;
   24380: out<=0;
   24381: out<=1;
   24382: out<=0;
   24383: out<=1;
   24384: out<=0;
   24385: out<=1;
   24386: out<=1;
   24387: out<=0;
   24388: out<=1;
   24389: out<=1;
   24390: out<=1;
   24391: out<=1;
   24392: out<=1;
   24393: out<=1;
   24394: out<=0;
   24395: out<=0;
   24396: out<=0;
   24397: out<=1;
   24398: out<=0;
   24399: out<=1;
   24400: out<=0;
   24401: out<=1;
   24402: out<=1;
   24403: out<=0;
   24404: out<=1;
   24405: out<=1;
   24406: out<=1;
   24407: out<=1;
   24408: out<=1;
   24409: out<=1;
   24410: out<=0;
   24411: out<=0;
   24412: out<=0;
   24413: out<=1;
   24414: out<=0;
   24415: out<=1;
   24416: out<=0;
   24417: out<=1;
   24418: out<=1;
   24419: out<=0;
   24420: out<=1;
   24421: out<=1;
   24422: out<=1;
   24423: out<=1;
   24424: out<=1;
   24425: out<=1;
   24426: out<=0;
   24427: out<=0;
   24428: out<=0;
   24429: out<=1;
   24430: out<=0;
   24431: out<=1;
   24432: out<=0;
   24433: out<=1;
   24434: out<=1;
   24435: out<=0;
   24436: out<=1;
   24437: out<=1;
   24438: out<=1;
   24439: out<=1;
   24440: out<=1;
   24441: out<=1;
   24442: out<=0;
   24443: out<=0;
   24444: out<=0;
   24445: out<=1;
   24446: out<=0;
   24447: out<=1;
   24448: out<=1;
   24449: out<=0;
   24450: out<=0;
   24451: out<=1;
   24452: out<=0;
   24453: out<=0;
   24454: out<=0;
   24455: out<=0;
   24456: out<=0;
   24457: out<=0;
   24458: out<=1;
   24459: out<=1;
   24460: out<=1;
   24461: out<=0;
   24462: out<=1;
   24463: out<=0;
   24464: out<=1;
   24465: out<=0;
   24466: out<=0;
   24467: out<=1;
   24468: out<=0;
   24469: out<=0;
   24470: out<=0;
   24471: out<=0;
   24472: out<=0;
   24473: out<=0;
   24474: out<=1;
   24475: out<=1;
   24476: out<=1;
   24477: out<=0;
   24478: out<=1;
   24479: out<=0;
   24480: out<=0;
   24481: out<=1;
   24482: out<=1;
   24483: out<=0;
   24484: out<=1;
   24485: out<=1;
   24486: out<=1;
   24487: out<=1;
   24488: out<=1;
   24489: out<=1;
   24490: out<=0;
   24491: out<=0;
   24492: out<=0;
   24493: out<=1;
   24494: out<=0;
   24495: out<=1;
   24496: out<=0;
   24497: out<=1;
   24498: out<=1;
   24499: out<=0;
   24500: out<=1;
   24501: out<=1;
   24502: out<=1;
   24503: out<=1;
   24504: out<=1;
   24505: out<=1;
   24506: out<=0;
   24507: out<=0;
   24508: out<=0;
   24509: out<=1;
   24510: out<=0;
   24511: out<=1;
   24512: out<=1;
   24513: out<=0;
   24514: out<=0;
   24515: out<=1;
   24516: out<=0;
   24517: out<=0;
   24518: out<=0;
   24519: out<=0;
   24520: out<=0;
   24521: out<=0;
   24522: out<=1;
   24523: out<=1;
   24524: out<=1;
   24525: out<=0;
   24526: out<=1;
   24527: out<=0;
   24528: out<=0;
   24529: out<=1;
   24530: out<=1;
   24531: out<=0;
   24532: out<=1;
   24533: out<=1;
   24534: out<=1;
   24535: out<=1;
   24536: out<=1;
   24537: out<=1;
   24538: out<=0;
   24539: out<=0;
   24540: out<=0;
   24541: out<=1;
   24542: out<=0;
   24543: out<=1;
   24544: out<=1;
   24545: out<=0;
   24546: out<=0;
   24547: out<=1;
   24548: out<=0;
   24549: out<=0;
   24550: out<=0;
   24551: out<=0;
   24552: out<=0;
   24553: out<=0;
   24554: out<=1;
   24555: out<=1;
   24556: out<=1;
   24557: out<=0;
   24558: out<=1;
   24559: out<=0;
   24560: out<=0;
   24561: out<=1;
   24562: out<=1;
   24563: out<=0;
   24564: out<=1;
   24565: out<=1;
   24566: out<=1;
   24567: out<=1;
   24568: out<=1;
   24569: out<=1;
   24570: out<=0;
   24571: out<=0;
   24572: out<=0;
   24573: out<=1;
   24574: out<=0;
   24575: out<=1;
   24576: out<=1;
   24577: out<=0;
   24578: out<=1;
   24579: out<=0;
   24580: out<=0;
   24581: out<=0;
   24582: out<=1;
   24583: out<=1;
   24584: out<=1;
   24585: out<=1;
   24586: out<=1;
   24587: out<=1;
   24588: out<=0;
   24589: out<=1;
   24590: out<=1;
   24591: out<=0;
   24592: out<=0;
   24593: out<=1;
   24594: out<=0;
   24595: out<=1;
   24596: out<=1;
   24597: out<=1;
   24598: out<=0;
   24599: out<=0;
   24600: out<=0;
   24601: out<=0;
   24602: out<=0;
   24603: out<=0;
   24604: out<=1;
   24605: out<=0;
   24606: out<=0;
   24607: out<=1;
   24608: out<=0;
   24609: out<=1;
   24610: out<=0;
   24611: out<=1;
   24612: out<=1;
   24613: out<=1;
   24614: out<=0;
   24615: out<=0;
   24616: out<=0;
   24617: out<=0;
   24618: out<=0;
   24619: out<=0;
   24620: out<=1;
   24621: out<=0;
   24622: out<=0;
   24623: out<=1;
   24624: out<=1;
   24625: out<=0;
   24626: out<=1;
   24627: out<=0;
   24628: out<=0;
   24629: out<=0;
   24630: out<=1;
   24631: out<=1;
   24632: out<=1;
   24633: out<=1;
   24634: out<=1;
   24635: out<=1;
   24636: out<=0;
   24637: out<=1;
   24638: out<=1;
   24639: out<=0;
   24640: out<=1;
   24641: out<=0;
   24642: out<=1;
   24643: out<=0;
   24644: out<=0;
   24645: out<=0;
   24646: out<=1;
   24647: out<=1;
   24648: out<=1;
   24649: out<=1;
   24650: out<=1;
   24651: out<=1;
   24652: out<=0;
   24653: out<=1;
   24654: out<=1;
   24655: out<=0;
   24656: out<=1;
   24657: out<=0;
   24658: out<=1;
   24659: out<=0;
   24660: out<=0;
   24661: out<=0;
   24662: out<=1;
   24663: out<=1;
   24664: out<=1;
   24665: out<=1;
   24666: out<=1;
   24667: out<=1;
   24668: out<=0;
   24669: out<=1;
   24670: out<=1;
   24671: out<=0;
   24672: out<=1;
   24673: out<=0;
   24674: out<=1;
   24675: out<=0;
   24676: out<=0;
   24677: out<=0;
   24678: out<=1;
   24679: out<=1;
   24680: out<=1;
   24681: out<=1;
   24682: out<=1;
   24683: out<=1;
   24684: out<=0;
   24685: out<=1;
   24686: out<=1;
   24687: out<=0;
   24688: out<=1;
   24689: out<=0;
   24690: out<=1;
   24691: out<=0;
   24692: out<=0;
   24693: out<=0;
   24694: out<=1;
   24695: out<=1;
   24696: out<=1;
   24697: out<=1;
   24698: out<=1;
   24699: out<=1;
   24700: out<=0;
   24701: out<=1;
   24702: out<=1;
   24703: out<=0;
   24704: out<=1;
   24705: out<=0;
   24706: out<=1;
   24707: out<=0;
   24708: out<=0;
   24709: out<=0;
   24710: out<=1;
   24711: out<=1;
   24712: out<=1;
   24713: out<=1;
   24714: out<=1;
   24715: out<=1;
   24716: out<=0;
   24717: out<=1;
   24718: out<=1;
   24719: out<=0;
   24720: out<=1;
   24721: out<=0;
   24722: out<=1;
   24723: out<=0;
   24724: out<=0;
   24725: out<=0;
   24726: out<=1;
   24727: out<=1;
   24728: out<=1;
   24729: out<=1;
   24730: out<=1;
   24731: out<=1;
   24732: out<=0;
   24733: out<=1;
   24734: out<=1;
   24735: out<=0;
   24736: out<=0;
   24737: out<=1;
   24738: out<=0;
   24739: out<=1;
   24740: out<=1;
   24741: out<=1;
   24742: out<=0;
   24743: out<=0;
   24744: out<=0;
   24745: out<=0;
   24746: out<=0;
   24747: out<=0;
   24748: out<=1;
   24749: out<=0;
   24750: out<=0;
   24751: out<=1;
   24752: out<=0;
   24753: out<=1;
   24754: out<=0;
   24755: out<=1;
   24756: out<=1;
   24757: out<=1;
   24758: out<=0;
   24759: out<=0;
   24760: out<=0;
   24761: out<=0;
   24762: out<=0;
   24763: out<=0;
   24764: out<=1;
   24765: out<=0;
   24766: out<=0;
   24767: out<=1;
   24768: out<=1;
   24769: out<=0;
   24770: out<=1;
   24771: out<=0;
   24772: out<=0;
   24773: out<=0;
   24774: out<=1;
   24775: out<=1;
   24776: out<=1;
   24777: out<=1;
   24778: out<=1;
   24779: out<=1;
   24780: out<=0;
   24781: out<=1;
   24782: out<=1;
   24783: out<=0;
   24784: out<=0;
   24785: out<=1;
   24786: out<=0;
   24787: out<=1;
   24788: out<=1;
   24789: out<=1;
   24790: out<=0;
   24791: out<=0;
   24792: out<=0;
   24793: out<=0;
   24794: out<=0;
   24795: out<=0;
   24796: out<=1;
   24797: out<=0;
   24798: out<=0;
   24799: out<=1;
   24800: out<=1;
   24801: out<=0;
   24802: out<=1;
   24803: out<=0;
   24804: out<=0;
   24805: out<=0;
   24806: out<=1;
   24807: out<=1;
   24808: out<=1;
   24809: out<=1;
   24810: out<=1;
   24811: out<=1;
   24812: out<=0;
   24813: out<=1;
   24814: out<=1;
   24815: out<=0;
   24816: out<=0;
   24817: out<=1;
   24818: out<=0;
   24819: out<=1;
   24820: out<=1;
   24821: out<=1;
   24822: out<=0;
   24823: out<=0;
   24824: out<=0;
   24825: out<=0;
   24826: out<=0;
   24827: out<=0;
   24828: out<=1;
   24829: out<=0;
   24830: out<=0;
   24831: out<=1;
   24832: out<=1;
   24833: out<=1;
   24834: out<=0;
   24835: out<=0;
   24836: out<=1;
   24837: out<=0;
   24838: out<=1;
   24839: out<=0;
   24840: out<=0;
   24841: out<=1;
   24842: out<=1;
   24843: out<=0;
   24844: out<=0;
   24845: out<=0;
   24846: out<=0;
   24847: out<=0;
   24848: out<=1;
   24849: out<=1;
   24850: out<=0;
   24851: out<=0;
   24852: out<=1;
   24853: out<=0;
   24854: out<=1;
   24855: out<=0;
   24856: out<=0;
   24857: out<=1;
   24858: out<=1;
   24859: out<=0;
   24860: out<=0;
   24861: out<=0;
   24862: out<=0;
   24863: out<=0;
   24864: out<=1;
   24865: out<=1;
   24866: out<=0;
   24867: out<=0;
   24868: out<=1;
   24869: out<=0;
   24870: out<=1;
   24871: out<=0;
   24872: out<=0;
   24873: out<=1;
   24874: out<=1;
   24875: out<=0;
   24876: out<=0;
   24877: out<=0;
   24878: out<=0;
   24879: out<=0;
   24880: out<=1;
   24881: out<=1;
   24882: out<=0;
   24883: out<=0;
   24884: out<=1;
   24885: out<=0;
   24886: out<=1;
   24887: out<=0;
   24888: out<=0;
   24889: out<=1;
   24890: out<=1;
   24891: out<=0;
   24892: out<=0;
   24893: out<=0;
   24894: out<=0;
   24895: out<=0;
   24896: out<=1;
   24897: out<=1;
   24898: out<=0;
   24899: out<=0;
   24900: out<=1;
   24901: out<=0;
   24902: out<=1;
   24903: out<=0;
   24904: out<=0;
   24905: out<=1;
   24906: out<=1;
   24907: out<=0;
   24908: out<=0;
   24909: out<=0;
   24910: out<=0;
   24911: out<=0;
   24912: out<=0;
   24913: out<=0;
   24914: out<=1;
   24915: out<=1;
   24916: out<=0;
   24917: out<=1;
   24918: out<=0;
   24919: out<=1;
   24920: out<=1;
   24921: out<=0;
   24922: out<=0;
   24923: out<=1;
   24924: out<=1;
   24925: out<=1;
   24926: out<=1;
   24927: out<=1;
   24928: out<=0;
   24929: out<=0;
   24930: out<=1;
   24931: out<=1;
   24932: out<=0;
   24933: out<=1;
   24934: out<=0;
   24935: out<=1;
   24936: out<=1;
   24937: out<=0;
   24938: out<=0;
   24939: out<=1;
   24940: out<=1;
   24941: out<=1;
   24942: out<=1;
   24943: out<=1;
   24944: out<=1;
   24945: out<=1;
   24946: out<=0;
   24947: out<=0;
   24948: out<=1;
   24949: out<=0;
   24950: out<=1;
   24951: out<=0;
   24952: out<=0;
   24953: out<=1;
   24954: out<=1;
   24955: out<=0;
   24956: out<=0;
   24957: out<=0;
   24958: out<=0;
   24959: out<=0;
   24960: out<=1;
   24961: out<=1;
   24962: out<=0;
   24963: out<=0;
   24964: out<=1;
   24965: out<=0;
   24966: out<=1;
   24967: out<=0;
   24968: out<=0;
   24969: out<=1;
   24970: out<=1;
   24971: out<=0;
   24972: out<=0;
   24973: out<=0;
   24974: out<=0;
   24975: out<=0;
   24976: out<=0;
   24977: out<=0;
   24978: out<=1;
   24979: out<=1;
   24980: out<=0;
   24981: out<=1;
   24982: out<=0;
   24983: out<=1;
   24984: out<=1;
   24985: out<=0;
   24986: out<=0;
   24987: out<=1;
   24988: out<=1;
   24989: out<=1;
   24990: out<=1;
   24991: out<=1;
   24992: out<=1;
   24993: out<=1;
   24994: out<=0;
   24995: out<=0;
   24996: out<=1;
   24997: out<=0;
   24998: out<=1;
   24999: out<=0;
   25000: out<=0;
   25001: out<=1;
   25002: out<=1;
   25003: out<=0;
   25004: out<=0;
   25005: out<=0;
   25006: out<=0;
   25007: out<=0;
   25008: out<=0;
   25009: out<=0;
   25010: out<=1;
   25011: out<=1;
   25012: out<=0;
   25013: out<=1;
   25014: out<=0;
   25015: out<=1;
   25016: out<=1;
   25017: out<=0;
   25018: out<=0;
   25019: out<=1;
   25020: out<=1;
   25021: out<=1;
   25022: out<=1;
   25023: out<=1;
   25024: out<=1;
   25025: out<=1;
   25026: out<=0;
   25027: out<=0;
   25028: out<=1;
   25029: out<=0;
   25030: out<=1;
   25031: out<=0;
   25032: out<=0;
   25033: out<=1;
   25034: out<=1;
   25035: out<=0;
   25036: out<=0;
   25037: out<=0;
   25038: out<=0;
   25039: out<=0;
   25040: out<=1;
   25041: out<=1;
   25042: out<=0;
   25043: out<=0;
   25044: out<=1;
   25045: out<=0;
   25046: out<=1;
   25047: out<=0;
   25048: out<=0;
   25049: out<=1;
   25050: out<=1;
   25051: out<=0;
   25052: out<=0;
   25053: out<=0;
   25054: out<=0;
   25055: out<=0;
   25056: out<=0;
   25057: out<=0;
   25058: out<=1;
   25059: out<=1;
   25060: out<=0;
   25061: out<=1;
   25062: out<=0;
   25063: out<=1;
   25064: out<=1;
   25065: out<=0;
   25066: out<=0;
   25067: out<=1;
   25068: out<=1;
   25069: out<=1;
   25070: out<=1;
   25071: out<=1;
   25072: out<=0;
   25073: out<=0;
   25074: out<=1;
   25075: out<=1;
   25076: out<=0;
   25077: out<=1;
   25078: out<=0;
   25079: out<=1;
   25080: out<=1;
   25081: out<=0;
   25082: out<=0;
   25083: out<=1;
   25084: out<=1;
   25085: out<=1;
   25086: out<=1;
   25087: out<=1;
   25088: out<=1;
   25089: out<=1;
   25090: out<=1;
   25091: out<=1;
   25092: out<=1;
   25093: out<=0;
   25094: out<=0;
   25095: out<=1;
   25096: out<=1;
   25097: out<=0;
   25098: out<=1;
   25099: out<=0;
   25100: out<=1;
   25101: out<=1;
   25102: out<=0;
   25103: out<=0;
   25104: out<=1;
   25105: out<=1;
   25106: out<=1;
   25107: out<=1;
   25108: out<=1;
   25109: out<=0;
   25110: out<=0;
   25111: out<=1;
   25112: out<=1;
   25113: out<=0;
   25114: out<=1;
   25115: out<=0;
   25116: out<=1;
   25117: out<=1;
   25118: out<=0;
   25119: out<=0;
   25120: out<=0;
   25121: out<=0;
   25122: out<=0;
   25123: out<=0;
   25124: out<=0;
   25125: out<=1;
   25126: out<=1;
   25127: out<=0;
   25128: out<=0;
   25129: out<=1;
   25130: out<=0;
   25131: out<=1;
   25132: out<=0;
   25133: out<=0;
   25134: out<=1;
   25135: out<=1;
   25136: out<=0;
   25137: out<=0;
   25138: out<=0;
   25139: out<=0;
   25140: out<=0;
   25141: out<=1;
   25142: out<=1;
   25143: out<=0;
   25144: out<=0;
   25145: out<=1;
   25146: out<=0;
   25147: out<=1;
   25148: out<=0;
   25149: out<=0;
   25150: out<=1;
   25151: out<=1;
   25152: out<=1;
   25153: out<=1;
   25154: out<=1;
   25155: out<=1;
   25156: out<=1;
   25157: out<=0;
   25158: out<=0;
   25159: out<=1;
   25160: out<=1;
   25161: out<=0;
   25162: out<=1;
   25163: out<=0;
   25164: out<=1;
   25165: out<=1;
   25166: out<=0;
   25167: out<=0;
   25168: out<=0;
   25169: out<=0;
   25170: out<=0;
   25171: out<=0;
   25172: out<=0;
   25173: out<=1;
   25174: out<=1;
   25175: out<=0;
   25176: out<=0;
   25177: out<=1;
   25178: out<=0;
   25179: out<=1;
   25180: out<=0;
   25181: out<=0;
   25182: out<=1;
   25183: out<=1;
   25184: out<=1;
   25185: out<=1;
   25186: out<=1;
   25187: out<=1;
   25188: out<=1;
   25189: out<=0;
   25190: out<=0;
   25191: out<=1;
   25192: out<=1;
   25193: out<=0;
   25194: out<=1;
   25195: out<=0;
   25196: out<=1;
   25197: out<=1;
   25198: out<=0;
   25199: out<=0;
   25200: out<=0;
   25201: out<=0;
   25202: out<=0;
   25203: out<=0;
   25204: out<=0;
   25205: out<=1;
   25206: out<=1;
   25207: out<=0;
   25208: out<=0;
   25209: out<=1;
   25210: out<=0;
   25211: out<=1;
   25212: out<=0;
   25213: out<=0;
   25214: out<=1;
   25215: out<=1;
   25216: out<=1;
   25217: out<=1;
   25218: out<=1;
   25219: out<=1;
   25220: out<=1;
   25221: out<=0;
   25222: out<=0;
   25223: out<=1;
   25224: out<=1;
   25225: out<=0;
   25226: out<=1;
   25227: out<=0;
   25228: out<=1;
   25229: out<=1;
   25230: out<=0;
   25231: out<=0;
   25232: out<=0;
   25233: out<=0;
   25234: out<=0;
   25235: out<=0;
   25236: out<=0;
   25237: out<=1;
   25238: out<=1;
   25239: out<=0;
   25240: out<=0;
   25241: out<=1;
   25242: out<=0;
   25243: out<=1;
   25244: out<=0;
   25245: out<=0;
   25246: out<=1;
   25247: out<=1;
   25248: out<=0;
   25249: out<=0;
   25250: out<=0;
   25251: out<=0;
   25252: out<=0;
   25253: out<=1;
   25254: out<=1;
   25255: out<=0;
   25256: out<=0;
   25257: out<=1;
   25258: out<=0;
   25259: out<=1;
   25260: out<=0;
   25261: out<=0;
   25262: out<=1;
   25263: out<=1;
   25264: out<=1;
   25265: out<=1;
   25266: out<=1;
   25267: out<=1;
   25268: out<=1;
   25269: out<=0;
   25270: out<=0;
   25271: out<=1;
   25272: out<=1;
   25273: out<=0;
   25274: out<=1;
   25275: out<=0;
   25276: out<=1;
   25277: out<=1;
   25278: out<=0;
   25279: out<=0;
   25280: out<=1;
   25281: out<=1;
   25282: out<=1;
   25283: out<=1;
   25284: out<=1;
   25285: out<=0;
   25286: out<=0;
   25287: out<=1;
   25288: out<=1;
   25289: out<=0;
   25290: out<=1;
   25291: out<=0;
   25292: out<=1;
   25293: out<=1;
   25294: out<=0;
   25295: out<=0;
   25296: out<=1;
   25297: out<=1;
   25298: out<=1;
   25299: out<=1;
   25300: out<=1;
   25301: out<=0;
   25302: out<=0;
   25303: out<=1;
   25304: out<=1;
   25305: out<=0;
   25306: out<=1;
   25307: out<=0;
   25308: out<=1;
   25309: out<=1;
   25310: out<=0;
   25311: out<=0;
   25312: out<=1;
   25313: out<=1;
   25314: out<=1;
   25315: out<=1;
   25316: out<=1;
   25317: out<=0;
   25318: out<=0;
   25319: out<=1;
   25320: out<=1;
   25321: out<=0;
   25322: out<=1;
   25323: out<=0;
   25324: out<=1;
   25325: out<=1;
   25326: out<=0;
   25327: out<=0;
   25328: out<=1;
   25329: out<=1;
   25330: out<=1;
   25331: out<=1;
   25332: out<=1;
   25333: out<=0;
   25334: out<=0;
   25335: out<=1;
   25336: out<=1;
   25337: out<=0;
   25338: out<=1;
   25339: out<=0;
   25340: out<=1;
   25341: out<=1;
   25342: out<=0;
   25343: out<=0;
   25344: out<=1;
   25345: out<=0;
   25346: out<=0;
   25347: out<=1;
   25348: out<=0;
   25349: out<=0;
   25350: out<=0;
   25351: out<=0;
   25352: out<=0;
   25353: out<=0;
   25354: out<=1;
   25355: out<=1;
   25356: out<=1;
   25357: out<=0;
   25358: out<=1;
   25359: out<=0;
   25360: out<=0;
   25361: out<=1;
   25362: out<=1;
   25363: out<=0;
   25364: out<=1;
   25365: out<=1;
   25366: out<=1;
   25367: out<=1;
   25368: out<=1;
   25369: out<=1;
   25370: out<=0;
   25371: out<=0;
   25372: out<=0;
   25373: out<=1;
   25374: out<=0;
   25375: out<=1;
   25376: out<=1;
   25377: out<=0;
   25378: out<=0;
   25379: out<=1;
   25380: out<=0;
   25381: out<=0;
   25382: out<=0;
   25383: out<=0;
   25384: out<=0;
   25385: out<=0;
   25386: out<=1;
   25387: out<=1;
   25388: out<=1;
   25389: out<=0;
   25390: out<=1;
   25391: out<=0;
   25392: out<=0;
   25393: out<=1;
   25394: out<=1;
   25395: out<=0;
   25396: out<=1;
   25397: out<=1;
   25398: out<=1;
   25399: out<=1;
   25400: out<=1;
   25401: out<=1;
   25402: out<=0;
   25403: out<=0;
   25404: out<=0;
   25405: out<=1;
   25406: out<=0;
   25407: out<=1;
   25408: out<=1;
   25409: out<=0;
   25410: out<=0;
   25411: out<=1;
   25412: out<=0;
   25413: out<=0;
   25414: out<=0;
   25415: out<=0;
   25416: out<=0;
   25417: out<=0;
   25418: out<=1;
   25419: out<=1;
   25420: out<=1;
   25421: out<=0;
   25422: out<=1;
   25423: out<=0;
   25424: out<=1;
   25425: out<=0;
   25426: out<=0;
   25427: out<=1;
   25428: out<=0;
   25429: out<=0;
   25430: out<=0;
   25431: out<=0;
   25432: out<=0;
   25433: out<=0;
   25434: out<=1;
   25435: out<=1;
   25436: out<=1;
   25437: out<=0;
   25438: out<=1;
   25439: out<=0;
   25440: out<=0;
   25441: out<=1;
   25442: out<=1;
   25443: out<=0;
   25444: out<=1;
   25445: out<=1;
   25446: out<=1;
   25447: out<=1;
   25448: out<=1;
   25449: out<=1;
   25450: out<=0;
   25451: out<=0;
   25452: out<=0;
   25453: out<=1;
   25454: out<=0;
   25455: out<=1;
   25456: out<=0;
   25457: out<=1;
   25458: out<=1;
   25459: out<=0;
   25460: out<=1;
   25461: out<=1;
   25462: out<=1;
   25463: out<=1;
   25464: out<=1;
   25465: out<=1;
   25466: out<=0;
   25467: out<=0;
   25468: out<=0;
   25469: out<=1;
   25470: out<=0;
   25471: out<=1;
   25472: out<=1;
   25473: out<=0;
   25474: out<=0;
   25475: out<=1;
   25476: out<=0;
   25477: out<=0;
   25478: out<=0;
   25479: out<=0;
   25480: out<=0;
   25481: out<=0;
   25482: out<=1;
   25483: out<=1;
   25484: out<=1;
   25485: out<=0;
   25486: out<=1;
   25487: out<=0;
   25488: out<=1;
   25489: out<=0;
   25490: out<=0;
   25491: out<=1;
   25492: out<=0;
   25493: out<=0;
   25494: out<=0;
   25495: out<=0;
   25496: out<=0;
   25497: out<=0;
   25498: out<=1;
   25499: out<=1;
   25500: out<=1;
   25501: out<=0;
   25502: out<=1;
   25503: out<=0;
   25504: out<=1;
   25505: out<=0;
   25506: out<=0;
   25507: out<=1;
   25508: out<=0;
   25509: out<=0;
   25510: out<=0;
   25511: out<=0;
   25512: out<=0;
   25513: out<=0;
   25514: out<=1;
   25515: out<=1;
   25516: out<=1;
   25517: out<=0;
   25518: out<=1;
   25519: out<=0;
   25520: out<=1;
   25521: out<=0;
   25522: out<=0;
   25523: out<=1;
   25524: out<=0;
   25525: out<=0;
   25526: out<=0;
   25527: out<=0;
   25528: out<=0;
   25529: out<=0;
   25530: out<=1;
   25531: out<=1;
   25532: out<=1;
   25533: out<=0;
   25534: out<=1;
   25535: out<=0;
   25536: out<=1;
   25537: out<=0;
   25538: out<=0;
   25539: out<=1;
   25540: out<=0;
   25541: out<=0;
   25542: out<=0;
   25543: out<=0;
   25544: out<=0;
   25545: out<=0;
   25546: out<=1;
   25547: out<=1;
   25548: out<=1;
   25549: out<=0;
   25550: out<=1;
   25551: out<=0;
   25552: out<=0;
   25553: out<=1;
   25554: out<=1;
   25555: out<=0;
   25556: out<=1;
   25557: out<=1;
   25558: out<=1;
   25559: out<=1;
   25560: out<=1;
   25561: out<=1;
   25562: out<=0;
   25563: out<=0;
   25564: out<=0;
   25565: out<=1;
   25566: out<=0;
   25567: out<=1;
   25568: out<=0;
   25569: out<=1;
   25570: out<=1;
   25571: out<=0;
   25572: out<=1;
   25573: out<=1;
   25574: out<=1;
   25575: out<=1;
   25576: out<=1;
   25577: out<=1;
   25578: out<=0;
   25579: out<=0;
   25580: out<=0;
   25581: out<=1;
   25582: out<=0;
   25583: out<=1;
   25584: out<=1;
   25585: out<=0;
   25586: out<=0;
   25587: out<=1;
   25588: out<=0;
   25589: out<=0;
   25590: out<=0;
   25591: out<=0;
   25592: out<=0;
   25593: out<=0;
   25594: out<=1;
   25595: out<=1;
   25596: out<=1;
   25597: out<=0;
   25598: out<=1;
   25599: out<=0;
   25600: out<=1;
   25601: out<=1;
   25602: out<=0;
   25603: out<=0;
   25604: out<=0;
   25605: out<=1;
   25606: out<=0;
   25607: out<=1;
   25608: out<=1;
   25609: out<=0;
   25610: out<=0;
   25611: out<=1;
   25612: out<=0;
   25613: out<=0;
   25614: out<=0;
   25615: out<=0;
   25616: out<=0;
   25617: out<=0;
   25618: out<=1;
   25619: out<=1;
   25620: out<=1;
   25621: out<=0;
   25622: out<=1;
   25623: out<=0;
   25624: out<=0;
   25625: out<=1;
   25626: out<=1;
   25627: out<=0;
   25628: out<=1;
   25629: out<=1;
   25630: out<=1;
   25631: out<=1;
   25632: out<=0;
   25633: out<=0;
   25634: out<=1;
   25635: out<=1;
   25636: out<=1;
   25637: out<=0;
   25638: out<=1;
   25639: out<=0;
   25640: out<=0;
   25641: out<=1;
   25642: out<=1;
   25643: out<=0;
   25644: out<=1;
   25645: out<=1;
   25646: out<=1;
   25647: out<=1;
   25648: out<=1;
   25649: out<=1;
   25650: out<=0;
   25651: out<=0;
   25652: out<=0;
   25653: out<=1;
   25654: out<=0;
   25655: out<=1;
   25656: out<=1;
   25657: out<=0;
   25658: out<=0;
   25659: out<=1;
   25660: out<=0;
   25661: out<=0;
   25662: out<=0;
   25663: out<=0;
   25664: out<=1;
   25665: out<=1;
   25666: out<=0;
   25667: out<=0;
   25668: out<=0;
   25669: out<=1;
   25670: out<=0;
   25671: out<=1;
   25672: out<=1;
   25673: out<=0;
   25674: out<=0;
   25675: out<=1;
   25676: out<=0;
   25677: out<=0;
   25678: out<=0;
   25679: out<=0;
   25680: out<=1;
   25681: out<=1;
   25682: out<=0;
   25683: out<=0;
   25684: out<=0;
   25685: out<=1;
   25686: out<=0;
   25687: out<=1;
   25688: out<=1;
   25689: out<=0;
   25690: out<=0;
   25691: out<=1;
   25692: out<=0;
   25693: out<=0;
   25694: out<=0;
   25695: out<=0;
   25696: out<=1;
   25697: out<=1;
   25698: out<=0;
   25699: out<=0;
   25700: out<=0;
   25701: out<=1;
   25702: out<=0;
   25703: out<=1;
   25704: out<=1;
   25705: out<=0;
   25706: out<=0;
   25707: out<=1;
   25708: out<=0;
   25709: out<=0;
   25710: out<=0;
   25711: out<=0;
   25712: out<=1;
   25713: out<=1;
   25714: out<=0;
   25715: out<=0;
   25716: out<=0;
   25717: out<=1;
   25718: out<=0;
   25719: out<=1;
   25720: out<=1;
   25721: out<=0;
   25722: out<=0;
   25723: out<=1;
   25724: out<=0;
   25725: out<=0;
   25726: out<=0;
   25727: out<=0;
   25728: out<=1;
   25729: out<=1;
   25730: out<=0;
   25731: out<=0;
   25732: out<=0;
   25733: out<=1;
   25734: out<=0;
   25735: out<=1;
   25736: out<=1;
   25737: out<=0;
   25738: out<=0;
   25739: out<=1;
   25740: out<=0;
   25741: out<=0;
   25742: out<=0;
   25743: out<=0;
   25744: out<=1;
   25745: out<=1;
   25746: out<=0;
   25747: out<=0;
   25748: out<=0;
   25749: out<=1;
   25750: out<=0;
   25751: out<=1;
   25752: out<=1;
   25753: out<=0;
   25754: out<=0;
   25755: out<=1;
   25756: out<=0;
   25757: out<=0;
   25758: out<=0;
   25759: out<=0;
   25760: out<=0;
   25761: out<=0;
   25762: out<=1;
   25763: out<=1;
   25764: out<=1;
   25765: out<=0;
   25766: out<=1;
   25767: out<=0;
   25768: out<=0;
   25769: out<=1;
   25770: out<=1;
   25771: out<=0;
   25772: out<=1;
   25773: out<=1;
   25774: out<=1;
   25775: out<=1;
   25776: out<=0;
   25777: out<=0;
   25778: out<=1;
   25779: out<=1;
   25780: out<=1;
   25781: out<=0;
   25782: out<=1;
   25783: out<=0;
   25784: out<=0;
   25785: out<=1;
   25786: out<=1;
   25787: out<=0;
   25788: out<=1;
   25789: out<=1;
   25790: out<=1;
   25791: out<=1;
   25792: out<=1;
   25793: out<=1;
   25794: out<=0;
   25795: out<=0;
   25796: out<=0;
   25797: out<=1;
   25798: out<=0;
   25799: out<=1;
   25800: out<=1;
   25801: out<=0;
   25802: out<=0;
   25803: out<=1;
   25804: out<=0;
   25805: out<=0;
   25806: out<=0;
   25807: out<=0;
   25808: out<=0;
   25809: out<=0;
   25810: out<=1;
   25811: out<=1;
   25812: out<=1;
   25813: out<=0;
   25814: out<=1;
   25815: out<=0;
   25816: out<=0;
   25817: out<=1;
   25818: out<=1;
   25819: out<=0;
   25820: out<=1;
   25821: out<=1;
   25822: out<=1;
   25823: out<=1;
   25824: out<=1;
   25825: out<=1;
   25826: out<=0;
   25827: out<=0;
   25828: out<=0;
   25829: out<=1;
   25830: out<=0;
   25831: out<=1;
   25832: out<=1;
   25833: out<=0;
   25834: out<=0;
   25835: out<=1;
   25836: out<=0;
   25837: out<=0;
   25838: out<=0;
   25839: out<=0;
   25840: out<=0;
   25841: out<=0;
   25842: out<=1;
   25843: out<=1;
   25844: out<=1;
   25845: out<=0;
   25846: out<=1;
   25847: out<=0;
   25848: out<=0;
   25849: out<=1;
   25850: out<=1;
   25851: out<=0;
   25852: out<=1;
   25853: out<=1;
   25854: out<=1;
   25855: out<=1;
   25856: out<=0;
   25857: out<=1;
   25858: out<=0;
   25859: out<=1;
   25860: out<=0;
   25861: out<=0;
   25862: out<=1;
   25863: out<=1;
   25864: out<=1;
   25865: out<=1;
   25866: out<=1;
   25867: out<=1;
   25868: out<=1;
   25869: out<=0;
   25870: out<=0;
   25871: out<=1;
   25872: out<=0;
   25873: out<=1;
   25874: out<=0;
   25875: out<=1;
   25876: out<=0;
   25877: out<=0;
   25878: out<=1;
   25879: out<=1;
   25880: out<=1;
   25881: out<=1;
   25882: out<=1;
   25883: out<=1;
   25884: out<=1;
   25885: out<=0;
   25886: out<=0;
   25887: out<=1;
   25888: out<=0;
   25889: out<=1;
   25890: out<=0;
   25891: out<=1;
   25892: out<=0;
   25893: out<=0;
   25894: out<=1;
   25895: out<=1;
   25896: out<=1;
   25897: out<=1;
   25898: out<=1;
   25899: out<=1;
   25900: out<=1;
   25901: out<=0;
   25902: out<=0;
   25903: out<=1;
   25904: out<=0;
   25905: out<=1;
   25906: out<=0;
   25907: out<=1;
   25908: out<=0;
   25909: out<=0;
   25910: out<=1;
   25911: out<=1;
   25912: out<=1;
   25913: out<=1;
   25914: out<=1;
   25915: out<=1;
   25916: out<=1;
   25917: out<=0;
   25918: out<=0;
   25919: out<=1;
   25920: out<=0;
   25921: out<=1;
   25922: out<=0;
   25923: out<=1;
   25924: out<=0;
   25925: out<=0;
   25926: out<=1;
   25927: out<=1;
   25928: out<=1;
   25929: out<=1;
   25930: out<=1;
   25931: out<=1;
   25932: out<=1;
   25933: out<=0;
   25934: out<=0;
   25935: out<=1;
   25936: out<=1;
   25937: out<=0;
   25938: out<=1;
   25939: out<=0;
   25940: out<=1;
   25941: out<=1;
   25942: out<=0;
   25943: out<=0;
   25944: out<=0;
   25945: out<=0;
   25946: out<=0;
   25947: out<=0;
   25948: out<=0;
   25949: out<=1;
   25950: out<=1;
   25951: out<=0;
   25952: out<=1;
   25953: out<=0;
   25954: out<=1;
   25955: out<=0;
   25956: out<=1;
   25957: out<=1;
   25958: out<=0;
   25959: out<=0;
   25960: out<=0;
   25961: out<=0;
   25962: out<=0;
   25963: out<=0;
   25964: out<=0;
   25965: out<=1;
   25966: out<=1;
   25967: out<=0;
   25968: out<=0;
   25969: out<=1;
   25970: out<=0;
   25971: out<=1;
   25972: out<=0;
   25973: out<=0;
   25974: out<=1;
   25975: out<=1;
   25976: out<=1;
   25977: out<=1;
   25978: out<=1;
   25979: out<=1;
   25980: out<=1;
   25981: out<=0;
   25982: out<=0;
   25983: out<=1;
   25984: out<=0;
   25985: out<=1;
   25986: out<=0;
   25987: out<=1;
   25988: out<=0;
   25989: out<=0;
   25990: out<=1;
   25991: out<=1;
   25992: out<=1;
   25993: out<=1;
   25994: out<=1;
   25995: out<=1;
   25996: out<=1;
   25997: out<=0;
   25998: out<=0;
   25999: out<=1;
   26000: out<=1;
   26001: out<=0;
   26002: out<=1;
   26003: out<=0;
   26004: out<=1;
   26005: out<=1;
   26006: out<=0;
   26007: out<=0;
   26008: out<=0;
   26009: out<=0;
   26010: out<=0;
   26011: out<=0;
   26012: out<=0;
   26013: out<=1;
   26014: out<=1;
   26015: out<=0;
   26016: out<=0;
   26017: out<=1;
   26018: out<=0;
   26019: out<=1;
   26020: out<=0;
   26021: out<=0;
   26022: out<=1;
   26023: out<=1;
   26024: out<=1;
   26025: out<=1;
   26026: out<=1;
   26027: out<=1;
   26028: out<=1;
   26029: out<=0;
   26030: out<=0;
   26031: out<=1;
   26032: out<=1;
   26033: out<=0;
   26034: out<=1;
   26035: out<=0;
   26036: out<=1;
   26037: out<=1;
   26038: out<=0;
   26039: out<=0;
   26040: out<=0;
   26041: out<=0;
   26042: out<=0;
   26043: out<=0;
   26044: out<=0;
   26045: out<=1;
   26046: out<=1;
   26047: out<=0;
   26048: out<=0;
   26049: out<=1;
   26050: out<=0;
   26051: out<=1;
   26052: out<=0;
   26053: out<=0;
   26054: out<=1;
   26055: out<=1;
   26056: out<=1;
   26057: out<=1;
   26058: out<=1;
   26059: out<=1;
   26060: out<=1;
   26061: out<=0;
   26062: out<=0;
   26063: out<=1;
   26064: out<=0;
   26065: out<=1;
   26066: out<=0;
   26067: out<=1;
   26068: out<=0;
   26069: out<=0;
   26070: out<=1;
   26071: out<=1;
   26072: out<=1;
   26073: out<=1;
   26074: out<=1;
   26075: out<=1;
   26076: out<=1;
   26077: out<=0;
   26078: out<=0;
   26079: out<=1;
   26080: out<=1;
   26081: out<=0;
   26082: out<=1;
   26083: out<=0;
   26084: out<=1;
   26085: out<=1;
   26086: out<=0;
   26087: out<=0;
   26088: out<=0;
   26089: out<=0;
   26090: out<=0;
   26091: out<=0;
   26092: out<=0;
   26093: out<=1;
   26094: out<=1;
   26095: out<=0;
   26096: out<=1;
   26097: out<=0;
   26098: out<=1;
   26099: out<=0;
   26100: out<=1;
   26101: out<=1;
   26102: out<=0;
   26103: out<=0;
   26104: out<=0;
   26105: out<=0;
   26106: out<=0;
   26107: out<=0;
   26108: out<=0;
   26109: out<=1;
   26110: out<=1;
   26111: out<=0;
   26112: out<=0;
   26113: out<=1;
   26114: out<=1;
   26115: out<=0;
   26116: out<=0;
   26117: out<=0;
   26118: out<=0;
   26119: out<=0;
   26120: out<=0;
   26121: out<=0;
   26122: out<=1;
   26123: out<=1;
   26124: out<=0;
   26125: out<=1;
   26126: out<=0;
   26127: out<=1;
   26128: out<=0;
   26129: out<=1;
   26130: out<=1;
   26131: out<=0;
   26132: out<=0;
   26133: out<=0;
   26134: out<=0;
   26135: out<=0;
   26136: out<=0;
   26137: out<=0;
   26138: out<=1;
   26139: out<=1;
   26140: out<=0;
   26141: out<=1;
   26142: out<=0;
   26143: out<=1;
   26144: out<=1;
   26145: out<=0;
   26146: out<=0;
   26147: out<=1;
   26148: out<=1;
   26149: out<=1;
   26150: out<=1;
   26151: out<=1;
   26152: out<=1;
   26153: out<=1;
   26154: out<=0;
   26155: out<=0;
   26156: out<=1;
   26157: out<=0;
   26158: out<=1;
   26159: out<=0;
   26160: out<=1;
   26161: out<=0;
   26162: out<=0;
   26163: out<=1;
   26164: out<=1;
   26165: out<=1;
   26166: out<=1;
   26167: out<=1;
   26168: out<=1;
   26169: out<=1;
   26170: out<=0;
   26171: out<=0;
   26172: out<=1;
   26173: out<=0;
   26174: out<=1;
   26175: out<=0;
   26176: out<=0;
   26177: out<=1;
   26178: out<=1;
   26179: out<=0;
   26180: out<=0;
   26181: out<=0;
   26182: out<=0;
   26183: out<=0;
   26184: out<=0;
   26185: out<=0;
   26186: out<=1;
   26187: out<=1;
   26188: out<=0;
   26189: out<=1;
   26190: out<=0;
   26191: out<=1;
   26192: out<=1;
   26193: out<=0;
   26194: out<=0;
   26195: out<=1;
   26196: out<=1;
   26197: out<=1;
   26198: out<=1;
   26199: out<=1;
   26200: out<=1;
   26201: out<=1;
   26202: out<=0;
   26203: out<=0;
   26204: out<=1;
   26205: out<=0;
   26206: out<=1;
   26207: out<=0;
   26208: out<=0;
   26209: out<=1;
   26210: out<=1;
   26211: out<=0;
   26212: out<=0;
   26213: out<=0;
   26214: out<=0;
   26215: out<=0;
   26216: out<=0;
   26217: out<=0;
   26218: out<=1;
   26219: out<=1;
   26220: out<=0;
   26221: out<=1;
   26222: out<=0;
   26223: out<=1;
   26224: out<=1;
   26225: out<=0;
   26226: out<=0;
   26227: out<=1;
   26228: out<=1;
   26229: out<=1;
   26230: out<=1;
   26231: out<=1;
   26232: out<=1;
   26233: out<=1;
   26234: out<=0;
   26235: out<=0;
   26236: out<=1;
   26237: out<=0;
   26238: out<=1;
   26239: out<=0;
   26240: out<=0;
   26241: out<=1;
   26242: out<=1;
   26243: out<=0;
   26244: out<=0;
   26245: out<=0;
   26246: out<=0;
   26247: out<=0;
   26248: out<=0;
   26249: out<=0;
   26250: out<=1;
   26251: out<=1;
   26252: out<=0;
   26253: out<=1;
   26254: out<=0;
   26255: out<=1;
   26256: out<=1;
   26257: out<=0;
   26258: out<=0;
   26259: out<=1;
   26260: out<=1;
   26261: out<=1;
   26262: out<=1;
   26263: out<=1;
   26264: out<=1;
   26265: out<=1;
   26266: out<=0;
   26267: out<=0;
   26268: out<=1;
   26269: out<=0;
   26270: out<=1;
   26271: out<=0;
   26272: out<=1;
   26273: out<=0;
   26274: out<=0;
   26275: out<=1;
   26276: out<=1;
   26277: out<=1;
   26278: out<=1;
   26279: out<=1;
   26280: out<=1;
   26281: out<=1;
   26282: out<=0;
   26283: out<=0;
   26284: out<=1;
   26285: out<=0;
   26286: out<=1;
   26287: out<=0;
   26288: out<=0;
   26289: out<=1;
   26290: out<=1;
   26291: out<=0;
   26292: out<=0;
   26293: out<=0;
   26294: out<=0;
   26295: out<=0;
   26296: out<=0;
   26297: out<=0;
   26298: out<=1;
   26299: out<=1;
   26300: out<=0;
   26301: out<=1;
   26302: out<=0;
   26303: out<=1;
   26304: out<=0;
   26305: out<=1;
   26306: out<=1;
   26307: out<=0;
   26308: out<=0;
   26309: out<=0;
   26310: out<=0;
   26311: out<=0;
   26312: out<=0;
   26313: out<=0;
   26314: out<=1;
   26315: out<=1;
   26316: out<=0;
   26317: out<=1;
   26318: out<=0;
   26319: out<=1;
   26320: out<=0;
   26321: out<=1;
   26322: out<=1;
   26323: out<=0;
   26324: out<=0;
   26325: out<=0;
   26326: out<=0;
   26327: out<=0;
   26328: out<=0;
   26329: out<=0;
   26330: out<=1;
   26331: out<=1;
   26332: out<=0;
   26333: out<=1;
   26334: out<=0;
   26335: out<=1;
   26336: out<=0;
   26337: out<=1;
   26338: out<=1;
   26339: out<=0;
   26340: out<=0;
   26341: out<=0;
   26342: out<=0;
   26343: out<=0;
   26344: out<=0;
   26345: out<=0;
   26346: out<=1;
   26347: out<=1;
   26348: out<=0;
   26349: out<=1;
   26350: out<=0;
   26351: out<=1;
   26352: out<=0;
   26353: out<=1;
   26354: out<=1;
   26355: out<=0;
   26356: out<=0;
   26357: out<=0;
   26358: out<=0;
   26359: out<=0;
   26360: out<=0;
   26361: out<=0;
   26362: out<=1;
   26363: out<=1;
   26364: out<=0;
   26365: out<=1;
   26366: out<=0;
   26367: out<=1;
   26368: out<=1;
   26369: out<=1;
   26370: out<=1;
   26371: out<=1;
   26372: out<=0;
   26373: out<=1;
   26374: out<=1;
   26375: out<=0;
   26376: out<=0;
   26377: out<=1;
   26378: out<=0;
   26379: out<=1;
   26380: out<=1;
   26381: out<=1;
   26382: out<=0;
   26383: out<=0;
   26384: out<=0;
   26385: out<=0;
   26386: out<=0;
   26387: out<=0;
   26388: out<=1;
   26389: out<=0;
   26390: out<=0;
   26391: out<=1;
   26392: out<=1;
   26393: out<=0;
   26394: out<=1;
   26395: out<=0;
   26396: out<=0;
   26397: out<=0;
   26398: out<=1;
   26399: out<=1;
   26400: out<=1;
   26401: out<=1;
   26402: out<=1;
   26403: out<=1;
   26404: out<=0;
   26405: out<=1;
   26406: out<=1;
   26407: out<=0;
   26408: out<=0;
   26409: out<=1;
   26410: out<=0;
   26411: out<=1;
   26412: out<=1;
   26413: out<=1;
   26414: out<=0;
   26415: out<=0;
   26416: out<=0;
   26417: out<=0;
   26418: out<=0;
   26419: out<=0;
   26420: out<=1;
   26421: out<=0;
   26422: out<=0;
   26423: out<=1;
   26424: out<=1;
   26425: out<=0;
   26426: out<=1;
   26427: out<=0;
   26428: out<=0;
   26429: out<=0;
   26430: out<=1;
   26431: out<=1;
   26432: out<=1;
   26433: out<=1;
   26434: out<=1;
   26435: out<=1;
   26436: out<=0;
   26437: out<=1;
   26438: out<=1;
   26439: out<=0;
   26440: out<=0;
   26441: out<=1;
   26442: out<=0;
   26443: out<=1;
   26444: out<=1;
   26445: out<=1;
   26446: out<=0;
   26447: out<=0;
   26448: out<=1;
   26449: out<=1;
   26450: out<=1;
   26451: out<=1;
   26452: out<=0;
   26453: out<=1;
   26454: out<=1;
   26455: out<=0;
   26456: out<=0;
   26457: out<=1;
   26458: out<=0;
   26459: out<=1;
   26460: out<=1;
   26461: out<=1;
   26462: out<=0;
   26463: out<=0;
   26464: out<=0;
   26465: out<=0;
   26466: out<=0;
   26467: out<=0;
   26468: out<=1;
   26469: out<=0;
   26470: out<=0;
   26471: out<=1;
   26472: out<=1;
   26473: out<=0;
   26474: out<=1;
   26475: out<=0;
   26476: out<=0;
   26477: out<=0;
   26478: out<=1;
   26479: out<=1;
   26480: out<=0;
   26481: out<=0;
   26482: out<=0;
   26483: out<=0;
   26484: out<=1;
   26485: out<=0;
   26486: out<=0;
   26487: out<=1;
   26488: out<=1;
   26489: out<=0;
   26490: out<=1;
   26491: out<=0;
   26492: out<=0;
   26493: out<=0;
   26494: out<=1;
   26495: out<=1;
   26496: out<=1;
   26497: out<=1;
   26498: out<=1;
   26499: out<=1;
   26500: out<=0;
   26501: out<=1;
   26502: out<=1;
   26503: out<=0;
   26504: out<=0;
   26505: out<=1;
   26506: out<=0;
   26507: out<=1;
   26508: out<=1;
   26509: out<=1;
   26510: out<=0;
   26511: out<=0;
   26512: out<=1;
   26513: out<=1;
   26514: out<=1;
   26515: out<=1;
   26516: out<=0;
   26517: out<=1;
   26518: out<=1;
   26519: out<=0;
   26520: out<=0;
   26521: out<=1;
   26522: out<=0;
   26523: out<=1;
   26524: out<=1;
   26525: out<=1;
   26526: out<=0;
   26527: out<=0;
   26528: out<=1;
   26529: out<=1;
   26530: out<=1;
   26531: out<=1;
   26532: out<=0;
   26533: out<=1;
   26534: out<=1;
   26535: out<=0;
   26536: out<=0;
   26537: out<=1;
   26538: out<=0;
   26539: out<=1;
   26540: out<=1;
   26541: out<=1;
   26542: out<=0;
   26543: out<=0;
   26544: out<=1;
   26545: out<=1;
   26546: out<=1;
   26547: out<=1;
   26548: out<=0;
   26549: out<=1;
   26550: out<=1;
   26551: out<=0;
   26552: out<=0;
   26553: out<=1;
   26554: out<=0;
   26555: out<=1;
   26556: out<=1;
   26557: out<=1;
   26558: out<=0;
   26559: out<=0;
   26560: out<=1;
   26561: out<=1;
   26562: out<=1;
   26563: out<=1;
   26564: out<=0;
   26565: out<=1;
   26566: out<=1;
   26567: out<=0;
   26568: out<=0;
   26569: out<=1;
   26570: out<=0;
   26571: out<=1;
   26572: out<=1;
   26573: out<=1;
   26574: out<=0;
   26575: out<=0;
   26576: out<=0;
   26577: out<=0;
   26578: out<=0;
   26579: out<=0;
   26580: out<=1;
   26581: out<=0;
   26582: out<=0;
   26583: out<=1;
   26584: out<=1;
   26585: out<=0;
   26586: out<=1;
   26587: out<=0;
   26588: out<=0;
   26589: out<=0;
   26590: out<=1;
   26591: out<=1;
   26592: out<=0;
   26593: out<=0;
   26594: out<=0;
   26595: out<=0;
   26596: out<=1;
   26597: out<=0;
   26598: out<=0;
   26599: out<=1;
   26600: out<=1;
   26601: out<=0;
   26602: out<=1;
   26603: out<=0;
   26604: out<=0;
   26605: out<=0;
   26606: out<=1;
   26607: out<=1;
   26608: out<=1;
   26609: out<=1;
   26610: out<=1;
   26611: out<=1;
   26612: out<=0;
   26613: out<=1;
   26614: out<=1;
   26615: out<=0;
   26616: out<=0;
   26617: out<=1;
   26618: out<=0;
   26619: out<=1;
   26620: out<=1;
   26621: out<=1;
   26622: out<=0;
   26623: out<=0;
   26624: out<=1;
   26625: out<=1;
   26626: out<=1;
   26627: out<=1;
   26628: out<=0;
   26629: out<=1;
   26630: out<=1;
   26631: out<=0;
   26632: out<=1;
   26633: out<=0;
   26634: out<=1;
   26635: out<=0;
   26636: out<=0;
   26637: out<=0;
   26638: out<=1;
   26639: out<=1;
   26640: out<=0;
   26641: out<=0;
   26642: out<=0;
   26643: out<=0;
   26644: out<=1;
   26645: out<=0;
   26646: out<=0;
   26647: out<=1;
   26648: out<=0;
   26649: out<=1;
   26650: out<=0;
   26651: out<=1;
   26652: out<=1;
   26653: out<=1;
   26654: out<=0;
   26655: out<=0;
   26656: out<=0;
   26657: out<=0;
   26658: out<=0;
   26659: out<=0;
   26660: out<=1;
   26661: out<=0;
   26662: out<=0;
   26663: out<=1;
   26664: out<=0;
   26665: out<=1;
   26666: out<=0;
   26667: out<=1;
   26668: out<=1;
   26669: out<=1;
   26670: out<=0;
   26671: out<=0;
   26672: out<=1;
   26673: out<=1;
   26674: out<=1;
   26675: out<=1;
   26676: out<=0;
   26677: out<=1;
   26678: out<=1;
   26679: out<=0;
   26680: out<=1;
   26681: out<=0;
   26682: out<=1;
   26683: out<=0;
   26684: out<=0;
   26685: out<=0;
   26686: out<=1;
   26687: out<=1;
   26688: out<=1;
   26689: out<=1;
   26690: out<=1;
   26691: out<=1;
   26692: out<=0;
   26693: out<=1;
   26694: out<=1;
   26695: out<=0;
   26696: out<=1;
   26697: out<=0;
   26698: out<=1;
   26699: out<=0;
   26700: out<=0;
   26701: out<=0;
   26702: out<=1;
   26703: out<=1;
   26704: out<=1;
   26705: out<=1;
   26706: out<=1;
   26707: out<=1;
   26708: out<=0;
   26709: out<=1;
   26710: out<=1;
   26711: out<=0;
   26712: out<=1;
   26713: out<=0;
   26714: out<=1;
   26715: out<=0;
   26716: out<=0;
   26717: out<=0;
   26718: out<=1;
   26719: out<=1;
   26720: out<=1;
   26721: out<=1;
   26722: out<=1;
   26723: out<=1;
   26724: out<=0;
   26725: out<=1;
   26726: out<=1;
   26727: out<=0;
   26728: out<=1;
   26729: out<=0;
   26730: out<=1;
   26731: out<=0;
   26732: out<=0;
   26733: out<=0;
   26734: out<=1;
   26735: out<=1;
   26736: out<=1;
   26737: out<=1;
   26738: out<=1;
   26739: out<=1;
   26740: out<=0;
   26741: out<=1;
   26742: out<=1;
   26743: out<=0;
   26744: out<=1;
   26745: out<=0;
   26746: out<=1;
   26747: out<=0;
   26748: out<=0;
   26749: out<=0;
   26750: out<=1;
   26751: out<=1;
   26752: out<=1;
   26753: out<=1;
   26754: out<=1;
   26755: out<=1;
   26756: out<=0;
   26757: out<=1;
   26758: out<=1;
   26759: out<=0;
   26760: out<=1;
   26761: out<=0;
   26762: out<=1;
   26763: out<=0;
   26764: out<=0;
   26765: out<=0;
   26766: out<=1;
   26767: out<=1;
   26768: out<=1;
   26769: out<=1;
   26770: out<=1;
   26771: out<=1;
   26772: out<=0;
   26773: out<=1;
   26774: out<=1;
   26775: out<=0;
   26776: out<=1;
   26777: out<=0;
   26778: out<=1;
   26779: out<=0;
   26780: out<=0;
   26781: out<=0;
   26782: out<=1;
   26783: out<=1;
   26784: out<=0;
   26785: out<=0;
   26786: out<=0;
   26787: out<=0;
   26788: out<=1;
   26789: out<=0;
   26790: out<=0;
   26791: out<=1;
   26792: out<=0;
   26793: out<=1;
   26794: out<=0;
   26795: out<=1;
   26796: out<=1;
   26797: out<=1;
   26798: out<=0;
   26799: out<=0;
   26800: out<=0;
   26801: out<=0;
   26802: out<=0;
   26803: out<=0;
   26804: out<=1;
   26805: out<=0;
   26806: out<=0;
   26807: out<=1;
   26808: out<=0;
   26809: out<=1;
   26810: out<=0;
   26811: out<=1;
   26812: out<=1;
   26813: out<=1;
   26814: out<=0;
   26815: out<=0;
   26816: out<=1;
   26817: out<=1;
   26818: out<=1;
   26819: out<=1;
   26820: out<=0;
   26821: out<=1;
   26822: out<=1;
   26823: out<=0;
   26824: out<=1;
   26825: out<=0;
   26826: out<=1;
   26827: out<=0;
   26828: out<=0;
   26829: out<=0;
   26830: out<=1;
   26831: out<=1;
   26832: out<=0;
   26833: out<=0;
   26834: out<=0;
   26835: out<=0;
   26836: out<=1;
   26837: out<=0;
   26838: out<=0;
   26839: out<=1;
   26840: out<=0;
   26841: out<=1;
   26842: out<=0;
   26843: out<=1;
   26844: out<=1;
   26845: out<=1;
   26846: out<=0;
   26847: out<=0;
   26848: out<=1;
   26849: out<=1;
   26850: out<=1;
   26851: out<=1;
   26852: out<=0;
   26853: out<=1;
   26854: out<=1;
   26855: out<=0;
   26856: out<=1;
   26857: out<=0;
   26858: out<=1;
   26859: out<=0;
   26860: out<=0;
   26861: out<=0;
   26862: out<=1;
   26863: out<=1;
   26864: out<=0;
   26865: out<=0;
   26866: out<=0;
   26867: out<=0;
   26868: out<=1;
   26869: out<=0;
   26870: out<=0;
   26871: out<=1;
   26872: out<=0;
   26873: out<=1;
   26874: out<=0;
   26875: out<=1;
   26876: out<=1;
   26877: out<=1;
   26878: out<=0;
   26879: out<=0;
   26880: out<=0;
   26881: out<=1;
   26882: out<=1;
   26883: out<=0;
   26884: out<=0;
   26885: out<=0;
   26886: out<=0;
   26887: out<=0;
   26888: out<=1;
   26889: out<=1;
   26890: out<=0;
   26891: out<=0;
   26892: out<=1;
   26893: out<=0;
   26894: out<=1;
   26895: out<=0;
   26896: out<=0;
   26897: out<=1;
   26898: out<=1;
   26899: out<=0;
   26900: out<=0;
   26901: out<=0;
   26902: out<=0;
   26903: out<=0;
   26904: out<=1;
   26905: out<=1;
   26906: out<=0;
   26907: out<=0;
   26908: out<=1;
   26909: out<=0;
   26910: out<=1;
   26911: out<=0;
   26912: out<=0;
   26913: out<=1;
   26914: out<=1;
   26915: out<=0;
   26916: out<=0;
   26917: out<=0;
   26918: out<=0;
   26919: out<=0;
   26920: out<=1;
   26921: out<=1;
   26922: out<=0;
   26923: out<=0;
   26924: out<=1;
   26925: out<=0;
   26926: out<=1;
   26927: out<=0;
   26928: out<=0;
   26929: out<=1;
   26930: out<=1;
   26931: out<=0;
   26932: out<=0;
   26933: out<=0;
   26934: out<=0;
   26935: out<=0;
   26936: out<=1;
   26937: out<=1;
   26938: out<=0;
   26939: out<=0;
   26940: out<=1;
   26941: out<=0;
   26942: out<=1;
   26943: out<=0;
   26944: out<=0;
   26945: out<=1;
   26946: out<=1;
   26947: out<=0;
   26948: out<=0;
   26949: out<=0;
   26950: out<=0;
   26951: out<=0;
   26952: out<=1;
   26953: out<=1;
   26954: out<=0;
   26955: out<=0;
   26956: out<=1;
   26957: out<=0;
   26958: out<=1;
   26959: out<=0;
   26960: out<=1;
   26961: out<=0;
   26962: out<=0;
   26963: out<=1;
   26964: out<=1;
   26965: out<=1;
   26966: out<=1;
   26967: out<=1;
   26968: out<=0;
   26969: out<=0;
   26970: out<=1;
   26971: out<=1;
   26972: out<=0;
   26973: out<=1;
   26974: out<=0;
   26975: out<=1;
   26976: out<=1;
   26977: out<=0;
   26978: out<=0;
   26979: out<=1;
   26980: out<=1;
   26981: out<=1;
   26982: out<=1;
   26983: out<=1;
   26984: out<=0;
   26985: out<=0;
   26986: out<=1;
   26987: out<=1;
   26988: out<=0;
   26989: out<=1;
   26990: out<=0;
   26991: out<=1;
   26992: out<=0;
   26993: out<=1;
   26994: out<=1;
   26995: out<=0;
   26996: out<=0;
   26997: out<=0;
   26998: out<=0;
   26999: out<=0;
   27000: out<=1;
   27001: out<=1;
   27002: out<=0;
   27003: out<=0;
   27004: out<=1;
   27005: out<=0;
   27006: out<=1;
   27007: out<=0;
   27008: out<=0;
   27009: out<=1;
   27010: out<=1;
   27011: out<=0;
   27012: out<=0;
   27013: out<=0;
   27014: out<=0;
   27015: out<=0;
   27016: out<=1;
   27017: out<=1;
   27018: out<=0;
   27019: out<=0;
   27020: out<=1;
   27021: out<=0;
   27022: out<=1;
   27023: out<=0;
   27024: out<=1;
   27025: out<=0;
   27026: out<=0;
   27027: out<=1;
   27028: out<=1;
   27029: out<=1;
   27030: out<=1;
   27031: out<=1;
   27032: out<=0;
   27033: out<=0;
   27034: out<=1;
   27035: out<=1;
   27036: out<=0;
   27037: out<=1;
   27038: out<=0;
   27039: out<=1;
   27040: out<=0;
   27041: out<=1;
   27042: out<=1;
   27043: out<=0;
   27044: out<=0;
   27045: out<=0;
   27046: out<=0;
   27047: out<=0;
   27048: out<=1;
   27049: out<=1;
   27050: out<=0;
   27051: out<=0;
   27052: out<=1;
   27053: out<=0;
   27054: out<=1;
   27055: out<=0;
   27056: out<=1;
   27057: out<=0;
   27058: out<=0;
   27059: out<=1;
   27060: out<=1;
   27061: out<=1;
   27062: out<=1;
   27063: out<=1;
   27064: out<=0;
   27065: out<=0;
   27066: out<=1;
   27067: out<=1;
   27068: out<=0;
   27069: out<=1;
   27070: out<=0;
   27071: out<=1;
   27072: out<=0;
   27073: out<=1;
   27074: out<=1;
   27075: out<=0;
   27076: out<=0;
   27077: out<=0;
   27078: out<=0;
   27079: out<=0;
   27080: out<=1;
   27081: out<=1;
   27082: out<=0;
   27083: out<=0;
   27084: out<=1;
   27085: out<=0;
   27086: out<=1;
   27087: out<=0;
   27088: out<=0;
   27089: out<=1;
   27090: out<=1;
   27091: out<=0;
   27092: out<=0;
   27093: out<=0;
   27094: out<=0;
   27095: out<=0;
   27096: out<=1;
   27097: out<=1;
   27098: out<=0;
   27099: out<=0;
   27100: out<=1;
   27101: out<=0;
   27102: out<=1;
   27103: out<=0;
   27104: out<=1;
   27105: out<=0;
   27106: out<=0;
   27107: out<=1;
   27108: out<=1;
   27109: out<=1;
   27110: out<=1;
   27111: out<=1;
   27112: out<=0;
   27113: out<=0;
   27114: out<=1;
   27115: out<=1;
   27116: out<=0;
   27117: out<=1;
   27118: out<=0;
   27119: out<=1;
   27120: out<=1;
   27121: out<=0;
   27122: out<=0;
   27123: out<=1;
   27124: out<=1;
   27125: out<=1;
   27126: out<=1;
   27127: out<=1;
   27128: out<=0;
   27129: out<=0;
   27130: out<=1;
   27131: out<=1;
   27132: out<=0;
   27133: out<=1;
   27134: out<=0;
   27135: out<=1;
   27136: out<=1;
   27137: out<=0;
   27138: out<=1;
   27139: out<=0;
   27140: out<=1;
   27141: out<=1;
   27142: out<=0;
   27143: out<=0;
   27144: out<=1;
   27145: out<=1;
   27146: out<=1;
   27147: out<=1;
   27148: out<=1;
   27149: out<=0;
   27150: out<=0;
   27151: out<=1;
   27152: out<=1;
   27153: out<=0;
   27154: out<=1;
   27155: out<=0;
   27156: out<=1;
   27157: out<=1;
   27158: out<=0;
   27159: out<=0;
   27160: out<=1;
   27161: out<=1;
   27162: out<=1;
   27163: out<=1;
   27164: out<=1;
   27165: out<=0;
   27166: out<=0;
   27167: out<=1;
   27168: out<=0;
   27169: out<=1;
   27170: out<=0;
   27171: out<=1;
   27172: out<=0;
   27173: out<=0;
   27174: out<=1;
   27175: out<=1;
   27176: out<=0;
   27177: out<=0;
   27178: out<=0;
   27179: out<=0;
   27180: out<=0;
   27181: out<=1;
   27182: out<=1;
   27183: out<=0;
   27184: out<=0;
   27185: out<=1;
   27186: out<=0;
   27187: out<=1;
   27188: out<=0;
   27189: out<=0;
   27190: out<=1;
   27191: out<=1;
   27192: out<=0;
   27193: out<=0;
   27194: out<=0;
   27195: out<=0;
   27196: out<=0;
   27197: out<=1;
   27198: out<=1;
   27199: out<=0;
   27200: out<=1;
   27201: out<=0;
   27202: out<=1;
   27203: out<=0;
   27204: out<=1;
   27205: out<=1;
   27206: out<=0;
   27207: out<=0;
   27208: out<=1;
   27209: out<=1;
   27210: out<=1;
   27211: out<=1;
   27212: out<=1;
   27213: out<=0;
   27214: out<=0;
   27215: out<=1;
   27216: out<=0;
   27217: out<=1;
   27218: out<=0;
   27219: out<=1;
   27220: out<=0;
   27221: out<=0;
   27222: out<=1;
   27223: out<=1;
   27224: out<=0;
   27225: out<=0;
   27226: out<=0;
   27227: out<=0;
   27228: out<=0;
   27229: out<=1;
   27230: out<=1;
   27231: out<=0;
   27232: out<=1;
   27233: out<=0;
   27234: out<=1;
   27235: out<=0;
   27236: out<=1;
   27237: out<=1;
   27238: out<=0;
   27239: out<=0;
   27240: out<=1;
   27241: out<=1;
   27242: out<=1;
   27243: out<=1;
   27244: out<=1;
   27245: out<=0;
   27246: out<=0;
   27247: out<=1;
   27248: out<=0;
   27249: out<=1;
   27250: out<=0;
   27251: out<=1;
   27252: out<=0;
   27253: out<=0;
   27254: out<=1;
   27255: out<=1;
   27256: out<=0;
   27257: out<=0;
   27258: out<=0;
   27259: out<=0;
   27260: out<=0;
   27261: out<=1;
   27262: out<=1;
   27263: out<=0;
   27264: out<=1;
   27265: out<=0;
   27266: out<=1;
   27267: out<=0;
   27268: out<=1;
   27269: out<=1;
   27270: out<=0;
   27271: out<=0;
   27272: out<=1;
   27273: out<=1;
   27274: out<=1;
   27275: out<=1;
   27276: out<=1;
   27277: out<=0;
   27278: out<=0;
   27279: out<=1;
   27280: out<=0;
   27281: out<=1;
   27282: out<=0;
   27283: out<=1;
   27284: out<=0;
   27285: out<=0;
   27286: out<=1;
   27287: out<=1;
   27288: out<=0;
   27289: out<=0;
   27290: out<=0;
   27291: out<=0;
   27292: out<=0;
   27293: out<=1;
   27294: out<=1;
   27295: out<=0;
   27296: out<=0;
   27297: out<=1;
   27298: out<=0;
   27299: out<=1;
   27300: out<=0;
   27301: out<=0;
   27302: out<=1;
   27303: out<=1;
   27304: out<=0;
   27305: out<=0;
   27306: out<=0;
   27307: out<=0;
   27308: out<=0;
   27309: out<=1;
   27310: out<=1;
   27311: out<=0;
   27312: out<=1;
   27313: out<=0;
   27314: out<=1;
   27315: out<=0;
   27316: out<=1;
   27317: out<=1;
   27318: out<=0;
   27319: out<=0;
   27320: out<=1;
   27321: out<=1;
   27322: out<=1;
   27323: out<=1;
   27324: out<=1;
   27325: out<=0;
   27326: out<=0;
   27327: out<=1;
   27328: out<=1;
   27329: out<=0;
   27330: out<=1;
   27331: out<=0;
   27332: out<=1;
   27333: out<=1;
   27334: out<=0;
   27335: out<=0;
   27336: out<=1;
   27337: out<=1;
   27338: out<=1;
   27339: out<=1;
   27340: out<=1;
   27341: out<=0;
   27342: out<=0;
   27343: out<=1;
   27344: out<=1;
   27345: out<=0;
   27346: out<=1;
   27347: out<=0;
   27348: out<=1;
   27349: out<=1;
   27350: out<=0;
   27351: out<=0;
   27352: out<=1;
   27353: out<=1;
   27354: out<=1;
   27355: out<=1;
   27356: out<=1;
   27357: out<=0;
   27358: out<=0;
   27359: out<=1;
   27360: out<=1;
   27361: out<=0;
   27362: out<=1;
   27363: out<=0;
   27364: out<=1;
   27365: out<=1;
   27366: out<=0;
   27367: out<=0;
   27368: out<=1;
   27369: out<=1;
   27370: out<=1;
   27371: out<=1;
   27372: out<=1;
   27373: out<=0;
   27374: out<=0;
   27375: out<=1;
   27376: out<=1;
   27377: out<=0;
   27378: out<=1;
   27379: out<=0;
   27380: out<=1;
   27381: out<=1;
   27382: out<=0;
   27383: out<=0;
   27384: out<=1;
   27385: out<=1;
   27386: out<=1;
   27387: out<=1;
   27388: out<=1;
   27389: out<=0;
   27390: out<=0;
   27391: out<=1;
   27392: out<=0;
   27393: out<=0;
   27394: out<=1;
   27395: out<=1;
   27396: out<=1;
   27397: out<=0;
   27398: out<=1;
   27399: out<=0;
   27400: out<=1;
   27401: out<=0;
   27402: out<=0;
   27403: out<=1;
   27404: out<=0;
   27405: out<=0;
   27406: out<=0;
   27407: out<=0;
   27408: out<=1;
   27409: out<=1;
   27410: out<=0;
   27411: out<=0;
   27412: out<=0;
   27413: out<=1;
   27414: out<=0;
   27415: out<=1;
   27416: out<=0;
   27417: out<=1;
   27418: out<=1;
   27419: out<=0;
   27420: out<=1;
   27421: out<=1;
   27422: out<=1;
   27423: out<=1;
   27424: out<=0;
   27425: out<=0;
   27426: out<=1;
   27427: out<=1;
   27428: out<=1;
   27429: out<=0;
   27430: out<=1;
   27431: out<=0;
   27432: out<=1;
   27433: out<=0;
   27434: out<=0;
   27435: out<=1;
   27436: out<=0;
   27437: out<=0;
   27438: out<=0;
   27439: out<=0;
   27440: out<=1;
   27441: out<=1;
   27442: out<=0;
   27443: out<=0;
   27444: out<=0;
   27445: out<=1;
   27446: out<=0;
   27447: out<=1;
   27448: out<=0;
   27449: out<=1;
   27450: out<=1;
   27451: out<=0;
   27452: out<=1;
   27453: out<=1;
   27454: out<=1;
   27455: out<=1;
   27456: out<=0;
   27457: out<=0;
   27458: out<=1;
   27459: out<=1;
   27460: out<=1;
   27461: out<=0;
   27462: out<=1;
   27463: out<=0;
   27464: out<=1;
   27465: out<=0;
   27466: out<=0;
   27467: out<=1;
   27468: out<=0;
   27469: out<=0;
   27470: out<=0;
   27471: out<=0;
   27472: out<=0;
   27473: out<=0;
   27474: out<=1;
   27475: out<=1;
   27476: out<=1;
   27477: out<=0;
   27478: out<=1;
   27479: out<=0;
   27480: out<=1;
   27481: out<=0;
   27482: out<=0;
   27483: out<=1;
   27484: out<=0;
   27485: out<=0;
   27486: out<=0;
   27487: out<=0;
   27488: out<=1;
   27489: out<=1;
   27490: out<=0;
   27491: out<=0;
   27492: out<=0;
   27493: out<=1;
   27494: out<=0;
   27495: out<=1;
   27496: out<=0;
   27497: out<=1;
   27498: out<=1;
   27499: out<=0;
   27500: out<=1;
   27501: out<=1;
   27502: out<=1;
   27503: out<=1;
   27504: out<=1;
   27505: out<=1;
   27506: out<=0;
   27507: out<=0;
   27508: out<=0;
   27509: out<=1;
   27510: out<=0;
   27511: out<=1;
   27512: out<=0;
   27513: out<=1;
   27514: out<=1;
   27515: out<=0;
   27516: out<=1;
   27517: out<=1;
   27518: out<=1;
   27519: out<=1;
   27520: out<=0;
   27521: out<=0;
   27522: out<=1;
   27523: out<=1;
   27524: out<=1;
   27525: out<=0;
   27526: out<=1;
   27527: out<=0;
   27528: out<=1;
   27529: out<=0;
   27530: out<=0;
   27531: out<=1;
   27532: out<=0;
   27533: out<=0;
   27534: out<=0;
   27535: out<=0;
   27536: out<=0;
   27537: out<=0;
   27538: out<=1;
   27539: out<=1;
   27540: out<=1;
   27541: out<=0;
   27542: out<=1;
   27543: out<=0;
   27544: out<=1;
   27545: out<=0;
   27546: out<=0;
   27547: out<=1;
   27548: out<=0;
   27549: out<=0;
   27550: out<=0;
   27551: out<=0;
   27552: out<=0;
   27553: out<=0;
   27554: out<=1;
   27555: out<=1;
   27556: out<=1;
   27557: out<=0;
   27558: out<=1;
   27559: out<=0;
   27560: out<=1;
   27561: out<=0;
   27562: out<=0;
   27563: out<=1;
   27564: out<=0;
   27565: out<=0;
   27566: out<=0;
   27567: out<=0;
   27568: out<=0;
   27569: out<=0;
   27570: out<=1;
   27571: out<=1;
   27572: out<=1;
   27573: out<=0;
   27574: out<=1;
   27575: out<=0;
   27576: out<=1;
   27577: out<=0;
   27578: out<=0;
   27579: out<=1;
   27580: out<=0;
   27581: out<=0;
   27582: out<=0;
   27583: out<=0;
   27584: out<=0;
   27585: out<=0;
   27586: out<=1;
   27587: out<=1;
   27588: out<=1;
   27589: out<=0;
   27590: out<=1;
   27591: out<=0;
   27592: out<=1;
   27593: out<=0;
   27594: out<=0;
   27595: out<=1;
   27596: out<=0;
   27597: out<=0;
   27598: out<=0;
   27599: out<=0;
   27600: out<=1;
   27601: out<=1;
   27602: out<=0;
   27603: out<=0;
   27604: out<=0;
   27605: out<=1;
   27606: out<=0;
   27607: out<=1;
   27608: out<=0;
   27609: out<=1;
   27610: out<=1;
   27611: out<=0;
   27612: out<=1;
   27613: out<=1;
   27614: out<=1;
   27615: out<=1;
   27616: out<=1;
   27617: out<=1;
   27618: out<=0;
   27619: out<=0;
   27620: out<=0;
   27621: out<=1;
   27622: out<=0;
   27623: out<=1;
   27624: out<=0;
   27625: out<=1;
   27626: out<=1;
   27627: out<=0;
   27628: out<=1;
   27629: out<=1;
   27630: out<=1;
   27631: out<=1;
   27632: out<=0;
   27633: out<=0;
   27634: out<=1;
   27635: out<=1;
   27636: out<=1;
   27637: out<=0;
   27638: out<=1;
   27639: out<=0;
   27640: out<=1;
   27641: out<=0;
   27642: out<=0;
   27643: out<=1;
   27644: out<=0;
   27645: out<=0;
   27646: out<=0;
   27647: out<=0;
   27648: out<=1;
   27649: out<=0;
   27650: out<=0;
   27651: out<=1;
   27652: out<=0;
   27653: out<=0;
   27654: out<=0;
   27655: out<=0;
   27656: out<=1;
   27657: out<=1;
   27658: out<=0;
   27659: out<=0;
   27660: out<=0;
   27661: out<=1;
   27662: out<=0;
   27663: out<=1;
   27664: out<=0;
   27665: out<=1;
   27666: out<=1;
   27667: out<=0;
   27668: out<=1;
   27669: out<=1;
   27670: out<=1;
   27671: out<=1;
   27672: out<=0;
   27673: out<=0;
   27674: out<=1;
   27675: out<=1;
   27676: out<=1;
   27677: out<=0;
   27678: out<=1;
   27679: out<=0;
   27680: out<=0;
   27681: out<=1;
   27682: out<=1;
   27683: out<=0;
   27684: out<=1;
   27685: out<=1;
   27686: out<=1;
   27687: out<=1;
   27688: out<=0;
   27689: out<=0;
   27690: out<=1;
   27691: out<=1;
   27692: out<=1;
   27693: out<=0;
   27694: out<=1;
   27695: out<=0;
   27696: out<=1;
   27697: out<=0;
   27698: out<=0;
   27699: out<=1;
   27700: out<=0;
   27701: out<=0;
   27702: out<=0;
   27703: out<=0;
   27704: out<=1;
   27705: out<=1;
   27706: out<=0;
   27707: out<=0;
   27708: out<=0;
   27709: out<=1;
   27710: out<=0;
   27711: out<=1;
   27712: out<=1;
   27713: out<=0;
   27714: out<=0;
   27715: out<=1;
   27716: out<=0;
   27717: out<=0;
   27718: out<=0;
   27719: out<=0;
   27720: out<=1;
   27721: out<=1;
   27722: out<=0;
   27723: out<=0;
   27724: out<=0;
   27725: out<=1;
   27726: out<=0;
   27727: out<=1;
   27728: out<=1;
   27729: out<=0;
   27730: out<=0;
   27731: out<=1;
   27732: out<=0;
   27733: out<=0;
   27734: out<=0;
   27735: out<=0;
   27736: out<=1;
   27737: out<=1;
   27738: out<=0;
   27739: out<=0;
   27740: out<=0;
   27741: out<=1;
   27742: out<=0;
   27743: out<=1;
   27744: out<=1;
   27745: out<=0;
   27746: out<=0;
   27747: out<=1;
   27748: out<=0;
   27749: out<=0;
   27750: out<=0;
   27751: out<=0;
   27752: out<=1;
   27753: out<=1;
   27754: out<=0;
   27755: out<=0;
   27756: out<=0;
   27757: out<=1;
   27758: out<=0;
   27759: out<=1;
   27760: out<=1;
   27761: out<=0;
   27762: out<=0;
   27763: out<=1;
   27764: out<=0;
   27765: out<=0;
   27766: out<=0;
   27767: out<=0;
   27768: out<=1;
   27769: out<=1;
   27770: out<=0;
   27771: out<=0;
   27772: out<=0;
   27773: out<=1;
   27774: out<=0;
   27775: out<=1;
   27776: out<=1;
   27777: out<=0;
   27778: out<=0;
   27779: out<=1;
   27780: out<=0;
   27781: out<=0;
   27782: out<=0;
   27783: out<=0;
   27784: out<=1;
   27785: out<=1;
   27786: out<=0;
   27787: out<=0;
   27788: out<=0;
   27789: out<=1;
   27790: out<=0;
   27791: out<=1;
   27792: out<=1;
   27793: out<=0;
   27794: out<=0;
   27795: out<=1;
   27796: out<=0;
   27797: out<=0;
   27798: out<=0;
   27799: out<=0;
   27800: out<=1;
   27801: out<=1;
   27802: out<=0;
   27803: out<=0;
   27804: out<=0;
   27805: out<=1;
   27806: out<=0;
   27807: out<=1;
   27808: out<=0;
   27809: out<=1;
   27810: out<=1;
   27811: out<=0;
   27812: out<=1;
   27813: out<=1;
   27814: out<=1;
   27815: out<=1;
   27816: out<=0;
   27817: out<=0;
   27818: out<=1;
   27819: out<=1;
   27820: out<=1;
   27821: out<=0;
   27822: out<=1;
   27823: out<=0;
   27824: out<=0;
   27825: out<=1;
   27826: out<=1;
   27827: out<=0;
   27828: out<=1;
   27829: out<=1;
   27830: out<=1;
   27831: out<=1;
   27832: out<=0;
   27833: out<=0;
   27834: out<=1;
   27835: out<=1;
   27836: out<=1;
   27837: out<=0;
   27838: out<=1;
   27839: out<=0;
   27840: out<=1;
   27841: out<=0;
   27842: out<=0;
   27843: out<=1;
   27844: out<=0;
   27845: out<=0;
   27846: out<=0;
   27847: out<=0;
   27848: out<=1;
   27849: out<=1;
   27850: out<=0;
   27851: out<=0;
   27852: out<=0;
   27853: out<=1;
   27854: out<=0;
   27855: out<=1;
   27856: out<=0;
   27857: out<=1;
   27858: out<=1;
   27859: out<=0;
   27860: out<=1;
   27861: out<=1;
   27862: out<=1;
   27863: out<=1;
   27864: out<=0;
   27865: out<=0;
   27866: out<=1;
   27867: out<=1;
   27868: out<=1;
   27869: out<=0;
   27870: out<=1;
   27871: out<=0;
   27872: out<=1;
   27873: out<=0;
   27874: out<=0;
   27875: out<=1;
   27876: out<=0;
   27877: out<=0;
   27878: out<=0;
   27879: out<=0;
   27880: out<=1;
   27881: out<=1;
   27882: out<=0;
   27883: out<=0;
   27884: out<=0;
   27885: out<=1;
   27886: out<=0;
   27887: out<=1;
   27888: out<=0;
   27889: out<=1;
   27890: out<=1;
   27891: out<=0;
   27892: out<=1;
   27893: out<=1;
   27894: out<=1;
   27895: out<=1;
   27896: out<=0;
   27897: out<=0;
   27898: out<=1;
   27899: out<=1;
   27900: out<=1;
   27901: out<=0;
   27902: out<=1;
   27903: out<=0;
   27904: out<=1;
   27905: out<=1;
   27906: out<=1;
   27907: out<=1;
   27908: out<=1;
   27909: out<=0;
   27910: out<=0;
   27911: out<=1;
   27912: out<=0;
   27913: out<=1;
   27914: out<=0;
   27915: out<=1;
   27916: out<=0;
   27917: out<=0;
   27918: out<=1;
   27919: out<=1;
   27920: out<=1;
   27921: out<=1;
   27922: out<=1;
   27923: out<=1;
   27924: out<=1;
   27925: out<=0;
   27926: out<=0;
   27927: out<=1;
   27928: out<=0;
   27929: out<=1;
   27930: out<=0;
   27931: out<=1;
   27932: out<=0;
   27933: out<=0;
   27934: out<=1;
   27935: out<=1;
   27936: out<=1;
   27937: out<=1;
   27938: out<=1;
   27939: out<=1;
   27940: out<=1;
   27941: out<=0;
   27942: out<=0;
   27943: out<=1;
   27944: out<=0;
   27945: out<=1;
   27946: out<=0;
   27947: out<=1;
   27948: out<=0;
   27949: out<=0;
   27950: out<=1;
   27951: out<=1;
   27952: out<=1;
   27953: out<=1;
   27954: out<=1;
   27955: out<=1;
   27956: out<=1;
   27957: out<=0;
   27958: out<=0;
   27959: out<=1;
   27960: out<=0;
   27961: out<=1;
   27962: out<=0;
   27963: out<=1;
   27964: out<=0;
   27965: out<=0;
   27966: out<=1;
   27967: out<=1;
   27968: out<=1;
   27969: out<=1;
   27970: out<=1;
   27971: out<=1;
   27972: out<=1;
   27973: out<=0;
   27974: out<=0;
   27975: out<=1;
   27976: out<=0;
   27977: out<=1;
   27978: out<=0;
   27979: out<=1;
   27980: out<=0;
   27981: out<=0;
   27982: out<=1;
   27983: out<=1;
   27984: out<=0;
   27985: out<=0;
   27986: out<=0;
   27987: out<=0;
   27988: out<=0;
   27989: out<=1;
   27990: out<=1;
   27991: out<=0;
   27992: out<=1;
   27993: out<=0;
   27994: out<=1;
   27995: out<=0;
   27996: out<=1;
   27997: out<=1;
   27998: out<=0;
   27999: out<=0;
   28000: out<=0;
   28001: out<=0;
   28002: out<=0;
   28003: out<=0;
   28004: out<=0;
   28005: out<=1;
   28006: out<=1;
   28007: out<=0;
   28008: out<=1;
   28009: out<=0;
   28010: out<=1;
   28011: out<=0;
   28012: out<=1;
   28013: out<=1;
   28014: out<=0;
   28015: out<=0;
   28016: out<=1;
   28017: out<=1;
   28018: out<=1;
   28019: out<=1;
   28020: out<=1;
   28021: out<=0;
   28022: out<=0;
   28023: out<=1;
   28024: out<=0;
   28025: out<=1;
   28026: out<=0;
   28027: out<=1;
   28028: out<=0;
   28029: out<=0;
   28030: out<=1;
   28031: out<=1;
   28032: out<=1;
   28033: out<=1;
   28034: out<=1;
   28035: out<=1;
   28036: out<=1;
   28037: out<=0;
   28038: out<=0;
   28039: out<=1;
   28040: out<=0;
   28041: out<=1;
   28042: out<=0;
   28043: out<=1;
   28044: out<=0;
   28045: out<=0;
   28046: out<=1;
   28047: out<=1;
   28048: out<=0;
   28049: out<=0;
   28050: out<=0;
   28051: out<=0;
   28052: out<=0;
   28053: out<=1;
   28054: out<=1;
   28055: out<=0;
   28056: out<=1;
   28057: out<=0;
   28058: out<=1;
   28059: out<=0;
   28060: out<=1;
   28061: out<=1;
   28062: out<=0;
   28063: out<=0;
   28064: out<=1;
   28065: out<=1;
   28066: out<=1;
   28067: out<=1;
   28068: out<=1;
   28069: out<=0;
   28070: out<=0;
   28071: out<=1;
   28072: out<=0;
   28073: out<=1;
   28074: out<=0;
   28075: out<=1;
   28076: out<=0;
   28077: out<=0;
   28078: out<=1;
   28079: out<=1;
   28080: out<=0;
   28081: out<=0;
   28082: out<=0;
   28083: out<=0;
   28084: out<=0;
   28085: out<=1;
   28086: out<=1;
   28087: out<=0;
   28088: out<=1;
   28089: out<=0;
   28090: out<=1;
   28091: out<=0;
   28092: out<=1;
   28093: out<=1;
   28094: out<=0;
   28095: out<=0;
   28096: out<=1;
   28097: out<=1;
   28098: out<=1;
   28099: out<=1;
   28100: out<=1;
   28101: out<=0;
   28102: out<=0;
   28103: out<=1;
   28104: out<=0;
   28105: out<=1;
   28106: out<=0;
   28107: out<=1;
   28108: out<=0;
   28109: out<=0;
   28110: out<=1;
   28111: out<=1;
   28112: out<=1;
   28113: out<=1;
   28114: out<=1;
   28115: out<=1;
   28116: out<=1;
   28117: out<=0;
   28118: out<=0;
   28119: out<=1;
   28120: out<=0;
   28121: out<=1;
   28122: out<=0;
   28123: out<=1;
   28124: out<=0;
   28125: out<=0;
   28126: out<=1;
   28127: out<=1;
   28128: out<=0;
   28129: out<=0;
   28130: out<=0;
   28131: out<=0;
   28132: out<=0;
   28133: out<=1;
   28134: out<=1;
   28135: out<=0;
   28136: out<=1;
   28137: out<=0;
   28138: out<=1;
   28139: out<=0;
   28140: out<=1;
   28141: out<=1;
   28142: out<=0;
   28143: out<=0;
   28144: out<=0;
   28145: out<=0;
   28146: out<=0;
   28147: out<=0;
   28148: out<=0;
   28149: out<=1;
   28150: out<=1;
   28151: out<=0;
   28152: out<=1;
   28153: out<=0;
   28154: out<=1;
   28155: out<=0;
   28156: out<=1;
   28157: out<=1;
   28158: out<=0;
   28159: out<=0;
   28160: out<=0;
   28161: out<=0;
   28162: out<=1;
   28163: out<=1;
   28164: out<=0;
   28165: out<=1;
   28166: out<=0;
   28167: out<=1;
   28168: out<=0;
   28169: out<=1;
   28170: out<=1;
   28171: out<=0;
   28172: out<=0;
   28173: out<=0;
   28174: out<=0;
   28175: out<=0;
   28176: out<=0;
   28177: out<=0;
   28178: out<=1;
   28179: out<=1;
   28180: out<=0;
   28181: out<=1;
   28182: out<=0;
   28183: out<=1;
   28184: out<=0;
   28185: out<=1;
   28186: out<=1;
   28187: out<=0;
   28188: out<=0;
   28189: out<=0;
   28190: out<=0;
   28191: out<=0;
   28192: out<=1;
   28193: out<=1;
   28194: out<=0;
   28195: out<=0;
   28196: out<=1;
   28197: out<=0;
   28198: out<=1;
   28199: out<=0;
   28200: out<=1;
   28201: out<=0;
   28202: out<=0;
   28203: out<=1;
   28204: out<=1;
   28205: out<=1;
   28206: out<=1;
   28207: out<=1;
   28208: out<=1;
   28209: out<=1;
   28210: out<=0;
   28211: out<=0;
   28212: out<=1;
   28213: out<=0;
   28214: out<=1;
   28215: out<=0;
   28216: out<=1;
   28217: out<=0;
   28218: out<=0;
   28219: out<=1;
   28220: out<=1;
   28221: out<=1;
   28222: out<=1;
   28223: out<=1;
   28224: out<=0;
   28225: out<=0;
   28226: out<=1;
   28227: out<=1;
   28228: out<=0;
   28229: out<=1;
   28230: out<=0;
   28231: out<=1;
   28232: out<=0;
   28233: out<=1;
   28234: out<=1;
   28235: out<=0;
   28236: out<=0;
   28237: out<=0;
   28238: out<=0;
   28239: out<=0;
   28240: out<=1;
   28241: out<=1;
   28242: out<=0;
   28243: out<=0;
   28244: out<=1;
   28245: out<=0;
   28246: out<=1;
   28247: out<=0;
   28248: out<=1;
   28249: out<=0;
   28250: out<=0;
   28251: out<=1;
   28252: out<=1;
   28253: out<=1;
   28254: out<=1;
   28255: out<=1;
   28256: out<=0;
   28257: out<=0;
   28258: out<=1;
   28259: out<=1;
   28260: out<=0;
   28261: out<=1;
   28262: out<=0;
   28263: out<=1;
   28264: out<=0;
   28265: out<=1;
   28266: out<=1;
   28267: out<=0;
   28268: out<=0;
   28269: out<=0;
   28270: out<=0;
   28271: out<=0;
   28272: out<=1;
   28273: out<=1;
   28274: out<=0;
   28275: out<=0;
   28276: out<=1;
   28277: out<=0;
   28278: out<=1;
   28279: out<=0;
   28280: out<=1;
   28281: out<=0;
   28282: out<=0;
   28283: out<=1;
   28284: out<=1;
   28285: out<=1;
   28286: out<=1;
   28287: out<=1;
   28288: out<=0;
   28289: out<=0;
   28290: out<=1;
   28291: out<=1;
   28292: out<=0;
   28293: out<=1;
   28294: out<=0;
   28295: out<=1;
   28296: out<=0;
   28297: out<=1;
   28298: out<=1;
   28299: out<=0;
   28300: out<=0;
   28301: out<=0;
   28302: out<=0;
   28303: out<=0;
   28304: out<=1;
   28305: out<=1;
   28306: out<=0;
   28307: out<=0;
   28308: out<=1;
   28309: out<=0;
   28310: out<=1;
   28311: out<=0;
   28312: out<=1;
   28313: out<=0;
   28314: out<=0;
   28315: out<=1;
   28316: out<=1;
   28317: out<=1;
   28318: out<=1;
   28319: out<=1;
   28320: out<=1;
   28321: out<=1;
   28322: out<=0;
   28323: out<=0;
   28324: out<=1;
   28325: out<=0;
   28326: out<=1;
   28327: out<=0;
   28328: out<=1;
   28329: out<=0;
   28330: out<=0;
   28331: out<=1;
   28332: out<=1;
   28333: out<=1;
   28334: out<=1;
   28335: out<=1;
   28336: out<=0;
   28337: out<=0;
   28338: out<=1;
   28339: out<=1;
   28340: out<=0;
   28341: out<=1;
   28342: out<=0;
   28343: out<=1;
   28344: out<=0;
   28345: out<=1;
   28346: out<=1;
   28347: out<=0;
   28348: out<=0;
   28349: out<=0;
   28350: out<=0;
   28351: out<=0;
   28352: out<=0;
   28353: out<=0;
   28354: out<=1;
   28355: out<=1;
   28356: out<=0;
   28357: out<=1;
   28358: out<=0;
   28359: out<=1;
   28360: out<=0;
   28361: out<=1;
   28362: out<=1;
   28363: out<=0;
   28364: out<=0;
   28365: out<=0;
   28366: out<=0;
   28367: out<=0;
   28368: out<=0;
   28369: out<=0;
   28370: out<=1;
   28371: out<=1;
   28372: out<=0;
   28373: out<=1;
   28374: out<=0;
   28375: out<=1;
   28376: out<=0;
   28377: out<=1;
   28378: out<=1;
   28379: out<=0;
   28380: out<=0;
   28381: out<=0;
   28382: out<=0;
   28383: out<=0;
   28384: out<=0;
   28385: out<=0;
   28386: out<=1;
   28387: out<=1;
   28388: out<=0;
   28389: out<=1;
   28390: out<=0;
   28391: out<=1;
   28392: out<=0;
   28393: out<=1;
   28394: out<=1;
   28395: out<=0;
   28396: out<=0;
   28397: out<=0;
   28398: out<=0;
   28399: out<=0;
   28400: out<=0;
   28401: out<=0;
   28402: out<=1;
   28403: out<=1;
   28404: out<=0;
   28405: out<=1;
   28406: out<=0;
   28407: out<=1;
   28408: out<=0;
   28409: out<=1;
   28410: out<=1;
   28411: out<=0;
   28412: out<=0;
   28413: out<=0;
   28414: out<=0;
   28415: out<=0;
   28416: out<=0;
   28417: out<=1;
   28418: out<=0;
   28419: out<=1;
   28420: out<=1;
   28421: out<=1;
   28422: out<=0;
   28423: out<=0;
   28424: out<=1;
   28425: out<=1;
   28426: out<=1;
   28427: out<=1;
   28428: out<=0;
   28429: out<=1;
   28430: out<=1;
   28431: out<=0;
   28432: out<=1;
   28433: out<=0;
   28434: out<=1;
   28435: out<=0;
   28436: out<=0;
   28437: out<=0;
   28438: out<=1;
   28439: out<=1;
   28440: out<=0;
   28441: out<=0;
   28442: out<=0;
   28443: out<=0;
   28444: out<=1;
   28445: out<=0;
   28446: out<=0;
   28447: out<=1;
   28448: out<=0;
   28449: out<=1;
   28450: out<=0;
   28451: out<=1;
   28452: out<=1;
   28453: out<=1;
   28454: out<=0;
   28455: out<=0;
   28456: out<=1;
   28457: out<=1;
   28458: out<=1;
   28459: out<=1;
   28460: out<=0;
   28461: out<=1;
   28462: out<=1;
   28463: out<=0;
   28464: out<=1;
   28465: out<=0;
   28466: out<=1;
   28467: out<=0;
   28468: out<=0;
   28469: out<=0;
   28470: out<=1;
   28471: out<=1;
   28472: out<=0;
   28473: out<=0;
   28474: out<=0;
   28475: out<=0;
   28476: out<=1;
   28477: out<=0;
   28478: out<=0;
   28479: out<=1;
   28480: out<=0;
   28481: out<=1;
   28482: out<=0;
   28483: out<=1;
   28484: out<=1;
   28485: out<=1;
   28486: out<=0;
   28487: out<=0;
   28488: out<=1;
   28489: out<=1;
   28490: out<=1;
   28491: out<=1;
   28492: out<=0;
   28493: out<=1;
   28494: out<=1;
   28495: out<=0;
   28496: out<=0;
   28497: out<=1;
   28498: out<=0;
   28499: out<=1;
   28500: out<=1;
   28501: out<=1;
   28502: out<=0;
   28503: out<=0;
   28504: out<=1;
   28505: out<=1;
   28506: out<=1;
   28507: out<=1;
   28508: out<=0;
   28509: out<=1;
   28510: out<=1;
   28511: out<=0;
   28512: out<=1;
   28513: out<=0;
   28514: out<=1;
   28515: out<=0;
   28516: out<=0;
   28517: out<=0;
   28518: out<=1;
   28519: out<=1;
   28520: out<=0;
   28521: out<=0;
   28522: out<=0;
   28523: out<=0;
   28524: out<=1;
   28525: out<=0;
   28526: out<=0;
   28527: out<=1;
   28528: out<=1;
   28529: out<=0;
   28530: out<=1;
   28531: out<=0;
   28532: out<=0;
   28533: out<=0;
   28534: out<=1;
   28535: out<=1;
   28536: out<=0;
   28537: out<=0;
   28538: out<=0;
   28539: out<=0;
   28540: out<=1;
   28541: out<=0;
   28542: out<=0;
   28543: out<=1;
   28544: out<=0;
   28545: out<=1;
   28546: out<=0;
   28547: out<=1;
   28548: out<=1;
   28549: out<=1;
   28550: out<=0;
   28551: out<=0;
   28552: out<=1;
   28553: out<=1;
   28554: out<=1;
   28555: out<=1;
   28556: out<=0;
   28557: out<=1;
   28558: out<=1;
   28559: out<=0;
   28560: out<=0;
   28561: out<=1;
   28562: out<=0;
   28563: out<=1;
   28564: out<=1;
   28565: out<=1;
   28566: out<=0;
   28567: out<=0;
   28568: out<=1;
   28569: out<=1;
   28570: out<=1;
   28571: out<=1;
   28572: out<=0;
   28573: out<=1;
   28574: out<=1;
   28575: out<=0;
   28576: out<=0;
   28577: out<=1;
   28578: out<=0;
   28579: out<=1;
   28580: out<=1;
   28581: out<=1;
   28582: out<=0;
   28583: out<=0;
   28584: out<=1;
   28585: out<=1;
   28586: out<=1;
   28587: out<=1;
   28588: out<=0;
   28589: out<=1;
   28590: out<=1;
   28591: out<=0;
   28592: out<=0;
   28593: out<=1;
   28594: out<=0;
   28595: out<=1;
   28596: out<=1;
   28597: out<=1;
   28598: out<=0;
   28599: out<=0;
   28600: out<=1;
   28601: out<=1;
   28602: out<=1;
   28603: out<=1;
   28604: out<=0;
   28605: out<=1;
   28606: out<=1;
   28607: out<=0;
   28608: out<=0;
   28609: out<=1;
   28610: out<=0;
   28611: out<=1;
   28612: out<=1;
   28613: out<=1;
   28614: out<=0;
   28615: out<=0;
   28616: out<=1;
   28617: out<=1;
   28618: out<=1;
   28619: out<=1;
   28620: out<=0;
   28621: out<=1;
   28622: out<=1;
   28623: out<=0;
   28624: out<=1;
   28625: out<=0;
   28626: out<=1;
   28627: out<=0;
   28628: out<=0;
   28629: out<=0;
   28630: out<=1;
   28631: out<=1;
   28632: out<=0;
   28633: out<=0;
   28634: out<=0;
   28635: out<=0;
   28636: out<=1;
   28637: out<=0;
   28638: out<=0;
   28639: out<=1;
   28640: out<=1;
   28641: out<=0;
   28642: out<=1;
   28643: out<=0;
   28644: out<=0;
   28645: out<=0;
   28646: out<=1;
   28647: out<=1;
   28648: out<=0;
   28649: out<=0;
   28650: out<=0;
   28651: out<=0;
   28652: out<=1;
   28653: out<=0;
   28654: out<=0;
   28655: out<=1;
   28656: out<=0;
   28657: out<=1;
   28658: out<=0;
   28659: out<=1;
   28660: out<=1;
   28661: out<=1;
   28662: out<=0;
   28663: out<=0;
   28664: out<=1;
   28665: out<=1;
   28666: out<=1;
   28667: out<=1;
   28668: out<=0;
   28669: out<=1;
   28670: out<=1;
   28671: out<=0;
   28672: out<=0;
   28673: out<=0;
   28674: out<=1;
   28675: out<=1;
   28676: out<=1;
   28677: out<=0;
   28678: out<=1;
   28679: out<=0;
   28680: out<=0;
   28681: out<=1;
   28682: out<=1;
   28683: out<=0;
   28684: out<=1;
   28685: out<=1;
   28686: out<=1;
   28687: out<=1;
   28688: out<=0;
   28689: out<=0;
   28690: out<=1;
   28691: out<=1;
   28692: out<=1;
   28693: out<=0;
   28694: out<=1;
   28695: out<=0;
   28696: out<=0;
   28697: out<=1;
   28698: out<=1;
   28699: out<=0;
   28700: out<=1;
   28701: out<=1;
   28702: out<=1;
   28703: out<=1;
   28704: out<=0;
   28705: out<=0;
   28706: out<=1;
   28707: out<=1;
   28708: out<=1;
   28709: out<=0;
   28710: out<=1;
   28711: out<=0;
   28712: out<=0;
   28713: out<=1;
   28714: out<=1;
   28715: out<=0;
   28716: out<=1;
   28717: out<=1;
   28718: out<=1;
   28719: out<=1;
   28720: out<=0;
   28721: out<=0;
   28722: out<=1;
   28723: out<=1;
   28724: out<=1;
   28725: out<=0;
   28726: out<=1;
   28727: out<=0;
   28728: out<=0;
   28729: out<=1;
   28730: out<=1;
   28731: out<=0;
   28732: out<=1;
   28733: out<=1;
   28734: out<=1;
   28735: out<=1;
   28736: out<=1;
   28737: out<=1;
   28738: out<=0;
   28739: out<=0;
   28740: out<=0;
   28741: out<=1;
   28742: out<=0;
   28743: out<=1;
   28744: out<=1;
   28745: out<=0;
   28746: out<=0;
   28747: out<=1;
   28748: out<=0;
   28749: out<=0;
   28750: out<=0;
   28751: out<=0;
   28752: out<=0;
   28753: out<=0;
   28754: out<=1;
   28755: out<=1;
   28756: out<=1;
   28757: out<=0;
   28758: out<=1;
   28759: out<=0;
   28760: out<=0;
   28761: out<=1;
   28762: out<=1;
   28763: out<=0;
   28764: out<=1;
   28765: out<=1;
   28766: out<=1;
   28767: out<=1;
   28768: out<=0;
   28769: out<=0;
   28770: out<=1;
   28771: out<=1;
   28772: out<=1;
   28773: out<=0;
   28774: out<=1;
   28775: out<=0;
   28776: out<=0;
   28777: out<=1;
   28778: out<=1;
   28779: out<=0;
   28780: out<=1;
   28781: out<=1;
   28782: out<=1;
   28783: out<=1;
   28784: out<=1;
   28785: out<=1;
   28786: out<=0;
   28787: out<=0;
   28788: out<=0;
   28789: out<=1;
   28790: out<=0;
   28791: out<=1;
   28792: out<=1;
   28793: out<=0;
   28794: out<=0;
   28795: out<=1;
   28796: out<=0;
   28797: out<=0;
   28798: out<=0;
   28799: out<=0;
   28800: out<=1;
   28801: out<=1;
   28802: out<=0;
   28803: out<=0;
   28804: out<=0;
   28805: out<=1;
   28806: out<=0;
   28807: out<=1;
   28808: out<=1;
   28809: out<=0;
   28810: out<=0;
   28811: out<=1;
   28812: out<=0;
   28813: out<=0;
   28814: out<=0;
   28815: out<=0;
   28816: out<=0;
   28817: out<=0;
   28818: out<=1;
   28819: out<=1;
   28820: out<=1;
   28821: out<=0;
   28822: out<=1;
   28823: out<=0;
   28824: out<=0;
   28825: out<=1;
   28826: out<=1;
   28827: out<=0;
   28828: out<=1;
   28829: out<=1;
   28830: out<=1;
   28831: out<=1;
   28832: out<=1;
   28833: out<=1;
   28834: out<=0;
   28835: out<=0;
   28836: out<=0;
   28837: out<=1;
   28838: out<=0;
   28839: out<=1;
   28840: out<=1;
   28841: out<=0;
   28842: out<=0;
   28843: out<=1;
   28844: out<=0;
   28845: out<=0;
   28846: out<=0;
   28847: out<=0;
   28848: out<=0;
   28849: out<=0;
   28850: out<=1;
   28851: out<=1;
   28852: out<=1;
   28853: out<=0;
   28854: out<=1;
   28855: out<=0;
   28856: out<=0;
   28857: out<=1;
   28858: out<=1;
   28859: out<=0;
   28860: out<=1;
   28861: out<=1;
   28862: out<=1;
   28863: out<=1;
   28864: out<=0;
   28865: out<=0;
   28866: out<=1;
   28867: out<=1;
   28868: out<=1;
   28869: out<=0;
   28870: out<=1;
   28871: out<=0;
   28872: out<=0;
   28873: out<=1;
   28874: out<=1;
   28875: out<=0;
   28876: out<=1;
   28877: out<=1;
   28878: out<=1;
   28879: out<=1;
   28880: out<=0;
   28881: out<=0;
   28882: out<=1;
   28883: out<=1;
   28884: out<=1;
   28885: out<=0;
   28886: out<=1;
   28887: out<=0;
   28888: out<=0;
   28889: out<=1;
   28890: out<=1;
   28891: out<=0;
   28892: out<=1;
   28893: out<=1;
   28894: out<=1;
   28895: out<=1;
   28896: out<=1;
   28897: out<=1;
   28898: out<=0;
   28899: out<=0;
   28900: out<=0;
   28901: out<=1;
   28902: out<=0;
   28903: out<=1;
   28904: out<=1;
   28905: out<=0;
   28906: out<=0;
   28907: out<=1;
   28908: out<=0;
   28909: out<=0;
   28910: out<=0;
   28911: out<=0;
   28912: out<=1;
   28913: out<=1;
   28914: out<=0;
   28915: out<=0;
   28916: out<=0;
   28917: out<=1;
   28918: out<=0;
   28919: out<=1;
   28920: out<=1;
   28921: out<=0;
   28922: out<=0;
   28923: out<=1;
   28924: out<=0;
   28925: out<=0;
   28926: out<=0;
   28927: out<=0;
   28928: out<=0;
   28929: out<=1;
   28930: out<=0;
   28931: out<=1;
   28932: out<=0;
   28933: out<=0;
   28934: out<=1;
   28935: out<=1;
   28936: out<=1;
   28937: out<=1;
   28938: out<=1;
   28939: out<=1;
   28940: out<=1;
   28941: out<=0;
   28942: out<=0;
   28943: out<=1;
   28944: out<=1;
   28945: out<=0;
   28946: out<=1;
   28947: out<=0;
   28948: out<=1;
   28949: out<=1;
   28950: out<=0;
   28951: out<=0;
   28952: out<=0;
   28953: out<=0;
   28954: out<=0;
   28955: out<=0;
   28956: out<=0;
   28957: out<=1;
   28958: out<=1;
   28959: out<=0;
   28960: out<=1;
   28961: out<=0;
   28962: out<=1;
   28963: out<=0;
   28964: out<=1;
   28965: out<=1;
   28966: out<=0;
   28967: out<=0;
   28968: out<=0;
   28969: out<=0;
   28970: out<=0;
   28971: out<=0;
   28972: out<=0;
   28973: out<=1;
   28974: out<=1;
   28975: out<=0;
   28976: out<=0;
   28977: out<=1;
   28978: out<=0;
   28979: out<=1;
   28980: out<=0;
   28981: out<=0;
   28982: out<=1;
   28983: out<=1;
   28984: out<=1;
   28985: out<=1;
   28986: out<=1;
   28987: out<=1;
   28988: out<=1;
   28989: out<=0;
   28990: out<=0;
   28991: out<=1;
   28992: out<=1;
   28993: out<=0;
   28994: out<=1;
   28995: out<=0;
   28996: out<=1;
   28997: out<=1;
   28998: out<=0;
   28999: out<=0;
   29000: out<=0;
   29001: out<=0;
   29002: out<=0;
   29003: out<=0;
   29004: out<=0;
   29005: out<=1;
   29006: out<=1;
   29007: out<=0;
   29008: out<=1;
   29009: out<=0;
   29010: out<=1;
   29011: out<=0;
   29012: out<=1;
   29013: out<=1;
   29014: out<=0;
   29015: out<=0;
   29016: out<=0;
   29017: out<=0;
   29018: out<=0;
   29019: out<=0;
   29020: out<=0;
   29021: out<=1;
   29022: out<=1;
   29023: out<=0;
   29024: out<=1;
   29025: out<=0;
   29026: out<=1;
   29027: out<=0;
   29028: out<=1;
   29029: out<=1;
   29030: out<=0;
   29031: out<=0;
   29032: out<=0;
   29033: out<=0;
   29034: out<=0;
   29035: out<=0;
   29036: out<=0;
   29037: out<=1;
   29038: out<=1;
   29039: out<=0;
   29040: out<=1;
   29041: out<=0;
   29042: out<=1;
   29043: out<=0;
   29044: out<=1;
   29045: out<=1;
   29046: out<=0;
   29047: out<=0;
   29048: out<=0;
   29049: out<=0;
   29050: out<=0;
   29051: out<=0;
   29052: out<=0;
   29053: out<=1;
   29054: out<=1;
   29055: out<=0;
   29056: out<=1;
   29057: out<=0;
   29058: out<=1;
   29059: out<=0;
   29060: out<=1;
   29061: out<=1;
   29062: out<=0;
   29063: out<=0;
   29064: out<=0;
   29065: out<=0;
   29066: out<=0;
   29067: out<=0;
   29068: out<=0;
   29069: out<=1;
   29070: out<=1;
   29071: out<=0;
   29072: out<=1;
   29073: out<=0;
   29074: out<=1;
   29075: out<=0;
   29076: out<=1;
   29077: out<=1;
   29078: out<=0;
   29079: out<=0;
   29080: out<=0;
   29081: out<=0;
   29082: out<=0;
   29083: out<=0;
   29084: out<=0;
   29085: out<=1;
   29086: out<=1;
   29087: out<=0;
   29088: out<=0;
   29089: out<=1;
   29090: out<=0;
   29091: out<=1;
   29092: out<=0;
   29093: out<=0;
   29094: out<=1;
   29095: out<=1;
   29096: out<=1;
   29097: out<=1;
   29098: out<=1;
   29099: out<=1;
   29100: out<=1;
   29101: out<=0;
   29102: out<=0;
   29103: out<=1;
   29104: out<=0;
   29105: out<=1;
   29106: out<=0;
   29107: out<=1;
   29108: out<=0;
   29109: out<=0;
   29110: out<=1;
   29111: out<=1;
   29112: out<=1;
   29113: out<=1;
   29114: out<=1;
   29115: out<=1;
   29116: out<=1;
   29117: out<=0;
   29118: out<=0;
   29119: out<=1;
   29120: out<=0;
   29121: out<=1;
   29122: out<=0;
   29123: out<=1;
   29124: out<=0;
   29125: out<=0;
   29126: out<=1;
   29127: out<=1;
   29128: out<=1;
   29129: out<=1;
   29130: out<=1;
   29131: out<=1;
   29132: out<=1;
   29133: out<=0;
   29134: out<=0;
   29135: out<=1;
   29136: out<=1;
   29137: out<=0;
   29138: out<=1;
   29139: out<=0;
   29140: out<=1;
   29141: out<=1;
   29142: out<=0;
   29143: out<=0;
   29144: out<=0;
   29145: out<=0;
   29146: out<=0;
   29147: out<=0;
   29148: out<=0;
   29149: out<=1;
   29150: out<=1;
   29151: out<=0;
   29152: out<=0;
   29153: out<=1;
   29154: out<=0;
   29155: out<=1;
   29156: out<=0;
   29157: out<=0;
   29158: out<=1;
   29159: out<=1;
   29160: out<=1;
   29161: out<=1;
   29162: out<=1;
   29163: out<=1;
   29164: out<=1;
   29165: out<=0;
   29166: out<=0;
   29167: out<=1;
   29168: out<=1;
   29169: out<=0;
   29170: out<=1;
   29171: out<=0;
   29172: out<=1;
   29173: out<=1;
   29174: out<=0;
   29175: out<=0;
   29176: out<=0;
   29177: out<=0;
   29178: out<=0;
   29179: out<=0;
   29180: out<=0;
   29181: out<=1;
   29182: out<=1;
   29183: out<=0;
   29184: out<=0;
   29185: out<=1;
   29186: out<=1;
   29187: out<=0;
   29188: out<=0;
   29189: out<=0;
   29190: out<=0;
   29191: out<=0;
   29192: out<=0;
   29193: out<=0;
   29194: out<=1;
   29195: out<=1;
   29196: out<=0;
   29197: out<=1;
   29198: out<=0;
   29199: out<=1;
   29200: out<=1;
   29201: out<=0;
   29202: out<=0;
   29203: out<=1;
   29204: out<=1;
   29205: out<=1;
   29206: out<=1;
   29207: out<=1;
   29208: out<=1;
   29209: out<=1;
   29210: out<=0;
   29211: out<=0;
   29212: out<=1;
   29213: out<=0;
   29214: out<=1;
   29215: out<=0;
   29216: out<=0;
   29217: out<=1;
   29218: out<=1;
   29219: out<=0;
   29220: out<=0;
   29221: out<=0;
   29222: out<=0;
   29223: out<=0;
   29224: out<=0;
   29225: out<=0;
   29226: out<=1;
   29227: out<=1;
   29228: out<=0;
   29229: out<=1;
   29230: out<=0;
   29231: out<=1;
   29232: out<=1;
   29233: out<=0;
   29234: out<=0;
   29235: out<=1;
   29236: out<=1;
   29237: out<=1;
   29238: out<=1;
   29239: out<=1;
   29240: out<=1;
   29241: out<=1;
   29242: out<=0;
   29243: out<=0;
   29244: out<=1;
   29245: out<=0;
   29246: out<=1;
   29247: out<=0;
   29248: out<=1;
   29249: out<=0;
   29250: out<=0;
   29251: out<=1;
   29252: out<=1;
   29253: out<=1;
   29254: out<=1;
   29255: out<=1;
   29256: out<=1;
   29257: out<=1;
   29258: out<=0;
   29259: out<=0;
   29260: out<=1;
   29261: out<=0;
   29262: out<=1;
   29263: out<=0;
   29264: out<=1;
   29265: out<=0;
   29266: out<=0;
   29267: out<=1;
   29268: out<=1;
   29269: out<=1;
   29270: out<=1;
   29271: out<=1;
   29272: out<=1;
   29273: out<=1;
   29274: out<=0;
   29275: out<=0;
   29276: out<=1;
   29277: out<=0;
   29278: out<=1;
   29279: out<=0;
   29280: out<=0;
   29281: out<=1;
   29282: out<=1;
   29283: out<=0;
   29284: out<=0;
   29285: out<=0;
   29286: out<=0;
   29287: out<=0;
   29288: out<=0;
   29289: out<=0;
   29290: out<=1;
   29291: out<=1;
   29292: out<=0;
   29293: out<=1;
   29294: out<=0;
   29295: out<=1;
   29296: out<=0;
   29297: out<=1;
   29298: out<=1;
   29299: out<=0;
   29300: out<=0;
   29301: out<=0;
   29302: out<=0;
   29303: out<=0;
   29304: out<=0;
   29305: out<=0;
   29306: out<=1;
   29307: out<=1;
   29308: out<=0;
   29309: out<=1;
   29310: out<=0;
   29311: out<=1;
   29312: out<=1;
   29313: out<=0;
   29314: out<=0;
   29315: out<=1;
   29316: out<=1;
   29317: out<=1;
   29318: out<=1;
   29319: out<=1;
   29320: out<=1;
   29321: out<=1;
   29322: out<=0;
   29323: out<=0;
   29324: out<=1;
   29325: out<=0;
   29326: out<=1;
   29327: out<=0;
   29328: out<=1;
   29329: out<=0;
   29330: out<=0;
   29331: out<=1;
   29332: out<=1;
   29333: out<=1;
   29334: out<=1;
   29335: out<=1;
   29336: out<=1;
   29337: out<=1;
   29338: out<=0;
   29339: out<=0;
   29340: out<=1;
   29341: out<=0;
   29342: out<=1;
   29343: out<=0;
   29344: out<=1;
   29345: out<=0;
   29346: out<=0;
   29347: out<=1;
   29348: out<=1;
   29349: out<=1;
   29350: out<=1;
   29351: out<=1;
   29352: out<=1;
   29353: out<=1;
   29354: out<=0;
   29355: out<=0;
   29356: out<=1;
   29357: out<=0;
   29358: out<=1;
   29359: out<=0;
   29360: out<=1;
   29361: out<=0;
   29362: out<=0;
   29363: out<=1;
   29364: out<=1;
   29365: out<=1;
   29366: out<=1;
   29367: out<=1;
   29368: out<=1;
   29369: out<=1;
   29370: out<=0;
   29371: out<=0;
   29372: out<=1;
   29373: out<=0;
   29374: out<=1;
   29375: out<=0;
   29376: out<=0;
   29377: out<=1;
   29378: out<=1;
   29379: out<=0;
   29380: out<=0;
   29381: out<=0;
   29382: out<=0;
   29383: out<=0;
   29384: out<=0;
   29385: out<=0;
   29386: out<=1;
   29387: out<=1;
   29388: out<=0;
   29389: out<=1;
   29390: out<=0;
   29391: out<=1;
   29392: out<=1;
   29393: out<=0;
   29394: out<=0;
   29395: out<=1;
   29396: out<=1;
   29397: out<=1;
   29398: out<=1;
   29399: out<=1;
   29400: out<=1;
   29401: out<=1;
   29402: out<=0;
   29403: out<=0;
   29404: out<=1;
   29405: out<=0;
   29406: out<=1;
   29407: out<=0;
   29408: out<=1;
   29409: out<=0;
   29410: out<=0;
   29411: out<=1;
   29412: out<=1;
   29413: out<=1;
   29414: out<=1;
   29415: out<=1;
   29416: out<=1;
   29417: out<=1;
   29418: out<=0;
   29419: out<=0;
   29420: out<=1;
   29421: out<=0;
   29422: out<=1;
   29423: out<=0;
   29424: out<=0;
   29425: out<=1;
   29426: out<=1;
   29427: out<=0;
   29428: out<=0;
   29429: out<=0;
   29430: out<=0;
   29431: out<=0;
   29432: out<=0;
   29433: out<=0;
   29434: out<=1;
   29435: out<=1;
   29436: out<=0;
   29437: out<=1;
   29438: out<=0;
   29439: out<=1;
   29440: out<=0;
   29441: out<=0;
   29442: out<=0;
   29443: out<=0;
   29444: out<=1;
   29445: out<=0;
   29446: out<=0;
   29447: out<=1;
   29448: out<=1;
   29449: out<=0;
   29450: out<=1;
   29451: out<=0;
   29452: out<=0;
   29453: out<=0;
   29454: out<=1;
   29455: out<=1;
   29456: out<=0;
   29457: out<=0;
   29458: out<=0;
   29459: out<=0;
   29460: out<=1;
   29461: out<=0;
   29462: out<=0;
   29463: out<=1;
   29464: out<=1;
   29465: out<=0;
   29466: out<=1;
   29467: out<=0;
   29468: out<=0;
   29469: out<=0;
   29470: out<=1;
   29471: out<=1;
   29472: out<=1;
   29473: out<=1;
   29474: out<=1;
   29475: out<=1;
   29476: out<=0;
   29477: out<=1;
   29478: out<=1;
   29479: out<=0;
   29480: out<=0;
   29481: out<=1;
   29482: out<=0;
   29483: out<=1;
   29484: out<=1;
   29485: out<=1;
   29486: out<=0;
   29487: out<=0;
   29488: out<=1;
   29489: out<=1;
   29490: out<=1;
   29491: out<=1;
   29492: out<=0;
   29493: out<=1;
   29494: out<=1;
   29495: out<=0;
   29496: out<=0;
   29497: out<=1;
   29498: out<=0;
   29499: out<=1;
   29500: out<=1;
   29501: out<=1;
   29502: out<=0;
   29503: out<=0;
   29504: out<=1;
   29505: out<=1;
   29506: out<=1;
   29507: out<=1;
   29508: out<=0;
   29509: out<=1;
   29510: out<=1;
   29511: out<=0;
   29512: out<=0;
   29513: out<=1;
   29514: out<=0;
   29515: out<=1;
   29516: out<=1;
   29517: out<=1;
   29518: out<=0;
   29519: out<=0;
   29520: out<=0;
   29521: out<=0;
   29522: out<=0;
   29523: out<=0;
   29524: out<=1;
   29525: out<=0;
   29526: out<=0;
   29527: out<=1;
   29528: out<=1;
   29529: out<=0;
   29530: out<=1;
   29531: out<=0;
   29532: out<=0;
   29533: out<=0;
   29534: out<=1;
   29535: out<=1;
   29536: out<=1;
   29537: out<=1;
   29538: out<=1;
   29539: out<=1;
   29540: out<=0;
   29541: out<=1;
   29542: out<=1;
   29543: out<=0;
   29544: out<=0;
   29545: out<=1;
   29546: out<=0;
   29547: out<=1;
   29548: out<=1;
   29549: out<=1;
   29550: out<=0;
   29551: out<=0;
   29552: out<=0;
   29553: out<=0;
   29554: out<=0;
   29555: out<=0;
   29556: out<=1;
   29557: out<=0;
   29558: out<=0;
   29559: out<=1;
   29560: out<=1;
   29561: out<=0;
   29562: out<=1;
   29563: out<=0;
   29564: out<=0;
   29565: out<=0;
   29566: out<=1;
   29567: out<=1;
   29568: out<=1;
   29569: out<=1;
   29570: out<=1;
   29571: out<=1;
   29572: out<=0;
   29573: out<=1;
   29574: out<=1;
   29575: out<=0;
   29576: out<=0;
   29577: out<=1;
   29578: out<=0;
   29579: out<=1;
   29580: out<=1;
   29581: out<=1;
   29582: out<=0;
   29583: out<=0;
   29584: out<=0;
   29585: out<=0;
   29586: out<=0;
   29587: out<=0;
   29588: out<=1;
   29589: out<=0;
   29590: out<=0;
   29591: out<=1;
   29592: out<=1;
   29593: out<=0;
   29594: out<=1;
   29595: out<=0;
   29596: out<=0;
   29597: out<=0;
   29598: out<=1;
   29599: out<=1;
   29600: out<=0;
   29601: out<=0;
   29602: out<=0;
   29603: out<=0;
   29604: out<=1;
   29605: out<=0;
   29606: out<=0;
   29607: out<=1;
   29608: out<=1;
   29609: out<=0;
   29610: out<=1;
   29611: out<=0;
   29612: out<=0;
   29613: out<=0;
   29614: out<=1;
   29615: out<=1;
   29616: out<=1;
   29617: out<=1;
   29618: out<=1;
   29619: out<=1;
   29620: out<=0;
   29621: out<=1;
   29622: out<=1;
   29623: out<=0;
   29624: out<=0;
   29625: out<=1;
   29626: out<=0;
   29627: out<=1;
   29628: out<=1;
   29629: out<=1;
   29630: out<=0;
   29631: out<=0;
   29632: out<=0;
   29633: out<=0;
   29634: out<=0;
   29635: out<=0;
   29636: out<=1;
   29637: out<=0;
   29638: out<=0;
   29639: out<=1;
   29640: out<=1;
   29641: out<=0;
   29642: out<=1;
   29643: out<=0;
   29644: out<=0;
   29645: out<=0;
   29646: out<=1;
   29647: out<=1;
   29648: out<=0;
   29649: out<=0;
   29650: out<=0;
   29651: out<=0;
   29652: out<=1;
   29653: out<=0;
   29654: out<=0;
   29655: out<=1;
   29656: out<=1;
   29657: out<=0;
   29658: out<=1;
   29659: out<=0;
   29660: out<=0;
   29661: out<=0;
   29662: out<=1;
   29663: out<=1;
   29664: out<=0;
   29665: out<=0;
   29666: out<=0;
   29667: out<=0;
   29668: out<=1;
   29669: out<=0;
   29670: out<=0;
   29671: out<=1;
   29672: out<=1;
   29673: out<=0;
   29674: out<=1;
   29675: out<=0;
   29676: out<=0;
   29677: out<=0;
   29678: out<=1;
   29679: out<=1;
   29680: out<=0;
   29681: out<=0;
   29682: out<=0;
   29683: out<=0;
   29684: out<=1;
   29685: out<=0;
   29686: out<=0;
   29687: out<=1;
   29688: out<=1;
   29689: out<=0;
   29690: out<=1;
   29691: out<=0;
   29692: out<=0;
   29693: out<=0;
   29694: out<=1;
   29695: out<=1;
   29696: out<=0;
   29697: out<=1;
   29698: out<=0;
   29699: out<=1;
   29700: out<=1;
   29701: out<=1;
   29702: out<=0;
   29703: out<=0;
   29704: out<=0;
   29705: out<=0;
   29706: out<=0;
   29707: out<=0;
   29708: out<=1;
   29709: out<=0;
   29710: out<=0;
   29711: out<=1;
   29712: out<=0;
   29713: out<=1;
   29714: out<=0;
   29715: out<=1;
   29716: out<=1;
   29717: out<=1;
   29718: out<=0;
   29719: out<=0;
   29720: out<=0;
   29721: out<=0;
   29722: out<=0;
   29723: out<=0;
   29724: out<=1;
   29725: out<=0;
   29726: out<=0;
   29727: out<=1;
   29728: out<=0;
   29729: out<=1;
   29730: out<=0;
   29731: out<=1;
   29732: out<=1;
   29733: out<=1;
   29734: out<=0;
   29735: out<=0;
   29736: out<=0;
   29737: out<=0;
   29738: out<=0;
   29739: out<=0;
   29740: out<=1;
   29741: out<=0;
   29742: out<=0;
   29743: out<=1;
   29744: out<=0;
   29745: out<=1;
   29746: out<=0;
   29747: out<=1;
   29748: out<=1;
   29749: out<=1;
   29750: out<=0;
   29751: out<=0;
   29752: out<=0;
   29753: out<=0;
   29754: out<=0;
   29755: out<=0;
   29756: out<=1;
   29757: out<=0;
   29758: out<=0;
   29759: out<=1;
   29760: out<=1;
   29761: out<=0;
   29762: out<=1;
   29763: out<=0;
   29764: out<=0;
   29765: out<=0;
   29766: out<=1;
   29767: out<=1;
   29768: out<=1;
   29769: out<=1;
   29770: out<=1;
   29771: out<=1;
   29772: out<=0;
   29773: out<=1;
   29774: out<=1;
   29775: out<=0;
   29776: out<=0;
   29777: out<=1;
   29778: out<=0;
   29779: out<=1;
   29780: out<=1;
   29781: out<=1;
   29782: out<=0;
   29783: out<=0;
   29784: out<=0;
   29785: out<=0;
   29786: out<=0;
   29787: out<=0;
   29788: out<=1;
   29789: out<=0;
   29790: out<=0;
   29791: out<=1;
   29792: out<=0;
   29793: out<=1;
   29794: out<=0;
   29795: out<=1;
   29796: out<=1;
   29797: out<=1;
   29798: out<=0;
   29799: out<=0;
   29800: out<=0;
   29801: out<=0;
   29802: out<=0;
   29803: out<=0;
   29804: out<=1;
   29805: out<=0;
   29806: out<=0;
   29807: out<=1;
   29808: out<=1;
   29809: out<=0;
   29810: out<=1;
   29811: out<=0;
   29812: out<=0;
   29813: out<=0;
   29814: out<=1;
   29815: out<=1;
   29816: out<=1;
   29817: out<=1;
   29818: out<=1;
   29819: out<=1;
   29820: out<=0;
   29821: out<=1;
   29822: out<=1;
   29823: out<=0;
   29824: out<=1;
   29825: out<=0;
   29826: out<=1;
   29827: out<=0;
   29828: out<=0;
   29829: out<=0;
   29830: out<=1;
   29831: out<=1;
   29832: out<=1;
   29833: out<=1;
   29834: out<=1;
   29835: out<=1;
   29836: out<=0;
   29837: out<=1;
   29838: out<=1;
   29839: out<=0;
   29840: out<=0;
   29841: out<=1;
   29842: out<=0;
   29843: out<=1;
   29844: out<=1;
   29845: out<=1;
   29846: out<=0;
   29847: out<=0;
   29848: out<=0;
   29849: out<=0;
   29850: out<=0;
   29851: out<=0;
   29852: out<=1;
   29853: out<=0;
   29854: out<=0;
   29855: out<=1;
   29856: out<=1;
   29857: out<=0;
   29858: out<=1;
   29859: out<=0;
   29860: out<=0;
   29861: out<=0;
   29862: out<=1;
   29863: out<=1;
   29864: out<=1;
   29865: out<=1;
   29866: out<=1;
   29867: out<=1;
   29868: out<=0;
   29869: out<=1;
   29870: out<=1;
   29871: out<=0;
   29872: out<=0;
   29873: out<=1;
   29874: out<=0;
   29875: out<=1;
   29876: out<=1;
   29877: out<=1;
   29878: out<=0;
   29879: out<=0;
   29880: out<=0;
   29881: out<=0;
   29882: out<=0;
   29883: out<=0;
   29884: out<=1;
   29885: out<=0;
   29886: out<=0;
   29887: out<=1;
   29888: out<=0;
   29889: out<=1;
   29890: out<=0;
   29891: out<=1;
   29892: out<=1;
   29893: out<=1;
   29894: out<=0;
   29895: out<=0;
   29896: out<=0;
   29897: out<=0;
   29898: out<=0;
   29899: out<=0;
   29900: out<=1;
   29901: out<=0;
   29902: out<=0;
   29903: out<=1;
   29904: out<=0;
   29905: out<=1;
   29906: out<=0;
   29907: out<=1;
   29908: out<=1;
   29909: out<=1;
   29910: out<=0;
   29911: out<=0;
   29912: out<=0;
   29913: out<=0;
   29914: out<=0;
   29915: out<=0;
   29916: out<=1;
   29917: out<=0;
   29918: out<=0;
   29919: out<=1;
   29920: out<=1;
   29921: out<=0;
   29922: out<=1;
   29923: out<=0;
   29924: out<=0;
   29925: out<=0;
   29926: out<=1;
   29927: out<=1;
   29928: out<=1;
   29929: out<=1;
   29930: out<=1;
   29931: out<=1;
   29932: out<=0;
   29933: out<=1;
   29934: out<=1;
   29935: out<=0;
   29936: out<=1;
   29937: out<=0;
   29938: out<=1;
   29939: out<=0;
   29940: out<=0;
   29941: out<=0;
   29942: out<=1;
   29943: out<=1;
   29944: out<=1;
   29945: out<=1;
   29946: out<=1;
   29947: out<=1;
   29948: out<=0;
   29949: out<=1;
   29950: out<=1;
   29951: out<=0;
   29952: out<=1;
   29953: out<=1;
   29954: out<=0;
   29955: out<=0;
   29956: out<=1;
   29957: out<=0;
   29958: out<=1;
   29959: out<=0;
   29960: out<=0;
   29961: out<=1;
   29962: out<=1;
   29963: out<=0;
   29964: out<=0;
   29965: out<=0;
   29966: out<=0;
   29967: out<=0;
   29968: out<=0;
   29969: out<=0;
   29970: out<=1;
   29971: out<=1;
   29972: out<=0;
   29973: out<=1;
   29974: out<=0;
   29975: out<=1;
   29976: out<=1;
   29977: out<=0;
   29978: out<=0;
   29979: out<=1;
   29980: out<=1;
   29981: out<=1;
   29982: out<=1;
   29983: out<=1;
   29984: out<=0;
   29985: out<=0;
   29986: out<=1;
   29987: out<=1;
   29988: out<=0;
   29989: out<=1;
   29990: out<=0;
   29991: out<=1;
   29992: out<=1;
   29993: out<=0;
   29994: out<=0;
   29995: out<=1;
   29996: out<=1;
   29997: out<=1;
   29998: out<=1;
   29999: out<=1;
   30000: out<=1;
   30001: out<=1;
   30002: out<=0;
   30003: out<=0;
   30004: out<=1;
   30005: out<=0;
   30006: out<=1;
   30007: out<=0;
   30008: out<=0;
   30009: out<=1;
   30010: out<=1;
   30011: out<=0;
   30012: out<=0;
   30013: out<=0;
   30014: out<=0;
   30015: out<=0;
   30016: out<=0;
   30017: out<=0;
   30018: out<=1;
   30019: out<=1;
   30020: out<=0;
   30021: out<=1;
   30022: out<=0;
   30023: out<=1;
   30024: out<=1;
   30025: out<=0;
   30026: out<=0;
   30027: out<=1;
   30028: out<=1;
   30029: out<=1;
   30030: out<=1;
   30031: out<=1;
   30032: out<=0;
   30033: out<=0;
   30034: out<=1;
   30035: out<=1;
   30036: out<=0;
   30037: out<=1;
   30038: out<=0;
   30039: out<=1;
   30040: out<=1;
   30041: out<=0;
   30042: out<=0;
   30043: out<=1;
   30044: out<=1;
   30045: out<=1;
   30046: out<=1;
   30047: out<=1;
   30048: out<=0;
   30049: out<=0;
   30050: out<=1;
   30051: out<=1;
   30052: out<=0;
   30053: out<=1;
   30054: out<=0;
   30055: out<=1;
   30056: out<=1;
   30057: out<=0;
   30058: out<=0;
   30059: out<=1;
   30060: out<=1;
   30061: out<=1;
   30062: out<=1;
   30063: out<=1;
   30064: out<=0;
   30065: out<=0;
   30066: out<=1;
   30067: out<=1;
   30068: out<=0;
   30069: out<=1;
   30070: out<=0;
   30071: out<=1;
   30072: out<=1;
   30073: out<=0;
   30074: out<=0;
   30075: out<=1;
   30076: out<=1;
   30077: out<=1;
   30078: out<=1;
   30079: out<=1;
   30080: out<=0;
   30081: out<=0;
   30082: out<=1;
   30083: out<=1;
   30084: out<=0;
   30085: out<=1;
   30086: out<=0;
   30087: out<=1;
   30088: out<=1;
   30089: out<=0;
   30090: out<=0;
   30091: out<=1;
   30092: out<=1;
   30093: out<=1;
   30094: out<=1;
   30095: out<=1;
   30096: out<=0;
   30097: out<=0;
   30098: out<=1;
   30099: out<=1;
   30100: out<=0;
   30101: out<=1;
   30102: out<=0;
   30103: out<=1;
   30104: out<=1;
   30105: out<=0;
   30106: out<=0;
   30107: out<=1;
   30108: out<=1;
   30109: out<=1;
   30110: out<=1;
   30111: out<=1;
   30112: out<=1;
   30113: out<=1;
   30114: out<=0;
   30115: out<=0;
   30116: out<=1;
   30117: out<=0;
   30118: out<=1;
   30119: out<=0;
   30120: out<=0;
   30121: out<=1;
   30122: out<=1;
   30123: out<=0;
   30124: out<=0;
   30125: out<=0;
   30126: out<=0;
   30127: out<=0;
   30128: out<=1;
   30129: out<=1;
   30130: out<=0;
   30131: out<=0;
   30132: out<=1;
   30133: out<=0;
   30134: out<=1;
   30135: out<=0;
   30136: out<=0;
   30137: out<=1;
   30138: out<=1;
   30139: out<=0;
   30140: out<=0;
   30141: out<=0;
   30142: out<=0;
   30143: out<=0;
   30144: out<=1;
   30145: out<=1;
   30146: out<=0;
   30147: out<=0;
   30148: out<=1;
   30149: out<=0;
   30150: out<=1;
   30151: out<=0;
   30152: out<=0;
   30153: out<=1;
   30154: out<=1;
   30155: out<=0;
   30156: out<=0;
   30157: out<=0;
   30158: out<=0;
   30159: out<=0;
   30160: out<=0;
   30161: out<=0;
   30162: out<=1;
   30163: out<=1;
   30164: out<=0;
   30165: out<=1;
   30166: out<=0;
   30167: out<=1;
   30168: out<=1;
   30169: out<=0;
   30170: out<=0;
   30171: out<=1;
   30172: out<=1;
   30173: out<=1;
   30174: out<=1;
   30175: out<=1;
   30176: out<=1;
   30177: out<=1;
   30178: out<=0;
   30179: out<=0;
   30180: out<=1;
   30181: out<=0;
   30182: out<=1;
   30183: out<=0;
   30184: out<=0;
   30185: out<=1;
   30186: out<=1;
   30187: out<=0;
   30188: out<=0;
   30189: out<=0;
   30190: out<=0;
   30191: out<=0;
   30192: out<=0;
   30193: out<=0;
   30194: out<=1;
   30195: out<=1;
   30196: out<=0;
   30197: out<=1;
   30198: out<=0;
   30199: out<=1;
   30200: out<=1;
   30201: out<=0;
   30202: out<=0;
   30203: out<=1;
   30204: out<=1;
   30205: out<=1;
   30206: out<=1;
   30207: out<=1;
   30208: out<=1;
   30209: out<=1;
   30210: out<=1;
   30211: out<=1;
   30212: out<=1;
   30213: out<=0;
   30214: out<=0;
   30215: out<=1;
   30216: out<=1;
   30217: out<=0;
   30218: out<=1;
   30219: out<=0;
   30220: out<=1;
   30221: out<=1;
   30222: out<=0;
   30223: out<=0;
   30224: out<=0;
   30225: out<=0;
   30226: out<=0;
   30227: out<=0;
   30228: out<=0;
   30229: out<=1;
   30230: out<=1;
   30231: out<=0;
   30232: out<=0;
   30233: out<=1;
   30234: out<=0;
   30235: out<=1;
   30236: out<=0;
   30237: out<=0;
   30238: out<=1;
   30239: out<=1;
   30240: out<=1;
   30241: out<=1;
   30242: out<=1;
   30243: out<=1;
   30244: out<=1;
   30245: out<=0;
   30246: out<=0;
   30247: out<=1;
   30248: out<=1;
   30249: out<=0;
   30250: out<=1;
   30251: out<=0;
   30252: out<=1;
   30253: out<=1;
   30254: out<=0;
   30255: out<=0;
   30256: out<=0;
   30257: out<=0;
   30258: out<=0;
   30259: out<=0;
   30260: out<=0;
   30261: out<=1;
   30262: out<=1;
   30263: out<=0;
   30264: out<=0;
   30265: out<=1;
   30266: out<=0;
   30267: out<=1;
   30268: out<=0;
   30269: out<=0;
   30270: out<=1;
   30271: out<=1;
   30272: out<=0;
   30273: out<=0;
   30274: out<=0;
   30275: out<=0;
   30276: out<=0;
   30277: out<=1;
   30278: out<=1;
   30279: out<=0;
   30280: out<=0;
   30281: out<=1;
   30282: out<=0;
   30283: out<=1;
   30284: out<=0;
   30285: out<=0;
   30286: out<=1;
   30287: out<=1;
   30288: out<=0;
   30289: out<=0;
   30290: out<=0;
   30291: out<=0;
   30292: out<=0;
   30293: out<=1;
   30294: out<=1;
   30295: out<=0;
   30296: out<=0;
   30297: out<=1;
   30298: out<=0;
   30299: out<=1;
   30300: out<=0;
   30301: out<=0;
   30302: out<=1;
   30303: out<=1;
   30304: out<=1;
   30305: out<=1;
   30306: out<=1;
   30307: out<=1;
   30308: out<=1;
   30309: out<=0;
   30310: out<=0;
   30311: out<=1;
   30312: out<=1;
   30313: out<=0;
   30314: out<=1;
   30315: out<=0;
   30316: out<=1;
   30317: out<=1;
   30318: out<=0;
   30319: out<=0;
   30320: out<=1;
   30321: out<=1;
   30322: out<=1;
   30323: out<=1;
   30324: out<=1;
   30325: out<=0;
   30326: out<=0;
   30327: out<=1;
   30328: out<=1;
   30329: out<=0;
   30330: out<=1;
   30331: out<=0;
   30332: out<=1;
   30333: out<=1;
   30334: out<=0;
   30335: out<=0;
   30336: out<=0;
   30337: out<=0;
   30338: out<=0;
   30339: out<=0;
   30340: out<=0;
   30341: out<=1;
   30342: out<=1;
   30343: out<=0;
   30344: out<=0;
   30345: out<=1;
   30346: out<=0;
   30347: out<=1;
   30348: out<=0;
   30349: out<=0;
   30350: out<=1;
   30351: out<=1;
   30352: out<=0;
   30353: out<=0;
   30354: out<=0;
   30355: out<=0;
   30356: out<=0;
   30357: out<=1;
   30358: out<=1;
   30359: out<=0;
   30360: out<=0;
   30361: out<=1;
   30362: out<=0;
   30363: out<=1;
   30364: out<=0;
   30365: out<=0;
   30366: out<=1;
   30367: out<=1;
   30368: out<=0;
   30369: out<=0;
   30370: out<=0;
   30371: out<=0;
   30372: out<=0;
   30373: out<=1;
   30374: out<=1;
   30375: out<=0;
   30376: out<=0;
   30377: out<=1;
   30378: out<=0;
   30379: out<=1;
   30380: out<=0;
   30381: out<=0;
   30382: out<=1;
   30383: out<=1;
   30384: out<=0;
   30385: out<=0;
   30386: out<=0;
   30387: out<=0;
   30388: out<=0;
   30389: out<=1;
   30390: out<=1;
   30391: out<=0;
   30392: out<=0;
   30393: out<=1;
   30394: out<=0;
   30395: out<=1;
   30396: out<=0;
   30397: out<=0;
   30398: out<=1;
   30399: out<=1;
   30400: out<=1;
   30401: out<=1;
   30402: out<=1;
   30403: out<=1;
   30404: out<=1;
   30405: out<=0;
   30406: out<=0;
   30407: out<=1;
   30408: out<=1;
   30409: out<=0;
   30410: out<=1;
   30411: out<=0;
   30412: out<=1;
   30413: out<=1;
   30414: out<=0;
   30415: out<=0;
   30416: out<=0;
   30417: out<=0;
   30418: out<=0;
   30419: out<=0;
   30420: out<=0;
   30421: out<=1;
   30422: out<=1;
   30423: out<=0;
   30424: out<=0;
   30425: out<=1;
   30426: out<=0;
   30427: out<=1;
   30428: out<=0;
   30429: out<=0;
   30430: out<=1;
   30431: out<=1;
   30432: out<=0;
   30433: out<=0;
   30434: out<=0;
   30435: out<=0;
   30436: out<=0;
   30437: out<=1;
   30438: out<=1;
   30439: out<=0;
   30440: out<=0;
   30441: out<=1;
   30442: out<=0;
   30443: out<=1;
   30444: out<=0;
   30445: out<=0;
   30446: out<=1;
   30447: out<=1;
   30448: out<=1;
   30449: out<=1;
   30450: out<=1;
   30451: out<=1;
   30452: out<=1;
   30453: out<=0;
   30454: out<=0;
   30455: out<=1;
   30456: out<=1;
   30457: out<=0;
   30458: out<=1;
   30459: out<=0;
   30460: out<=1;
   30461: out<=1;
   30462: out<=0;
   30463: out<=0;
   30464: out<=0;
   30465: out<=1;
   30466: out<=1;
   30467: out<=0;
   30468: out<=1;
   30469: out<=1;
   30470: out<=1;
   30471: out<=1;
   30472: out<=1;
   30473: out<=1;
   30474: out<=0;
   30475: out<=0;
   30476: out<=0;
   30477: out<=1;
   30478: out<=0;
   30479: out<=1;
   30480: out<=0;
   30481: out<=1;
   30482: out<=1;
   30483: out<=0;
   30484: out<=1;
   30485: out<=1;
   30486: out<=1;
   30487: out<=1;
   30488: out<=1;
   30489: out<=1;
   30490: out<=0;
   30491: out<=0;
   30492: out<=0;
   30493: out<=1;
   30494: out<=0;
   30495: out<=1;
   30496: out<=1;
   30497: out<=0;
   30498: out<=0;
   30499: out<=1;
   30500: out<=0;
   30501: out<=0;
   30502: out<=0;
   30503: out<=0;
   30504: out<=0;
   30505: out<=0;
   30506: out<=1;
   30507: out<=1;
   30508: out<=1;
   30509: out<=0;
   30510: out<=1;
   30511: out<=0;
   30512: out<=1;
   30513: out<=0;
   30514: out<=0;
   30515: out<=1;
   30516: out<=0;
   30517: out<=0;
   30518: out<=0;
   30519: out<=0;
   30520: out<=0;
   30521: out<=0;
   30522: out<=1;
   30523: out<=1;
   30524: out<=1;
   30525: out<=0;
   30526: out<=1;
   30527: out<=0;
   30528: out<=1;
   30529: out<=0;
   30530: out<=0;
   30531: out<=1;
   30532: out<=0;
   30533: out<=0;
   30534: out<=0;
   30535: out<=0;
   30536: out<=0;
   30537: out<=0;
   30538: out<=1;
   30539: out<=1;
   30540: out<=1;
   30541: out<=0;
   30542: out<=1;
   30543: out<=0;
   30544: out<=0;
   30545: out<=1;
   30546: out<=1;
   30547: out<=0;
   30548: out<=1;
   30549: out<=1;
   30550: out<=1;
   30551: out<=1;
   30552: out<=1;
   30553: out<=1;
   30554: out<=0;
   30555: out<=0;
   30556: out<=0;
   30557: out<=1;
   30558: out<=0;
   30559: out<=1;
   30560: out<=1;
   30561: out<=0;
   30562: out<=0;
   30563: out<=1;
   30564: out<=0;
   30565: out<=0;
   30566: out<=0;
   30567: out<=0;
   30568: out<=0;
   30569: out<=0;
   30570: out<=1;
   30571: out<=1;
   30572: out<=1;
   30573: out<=0;
   30574: out<=1;
   30575: out<=0;
   30576: out<=0;
   30577: out<=1;
   30578: out<=1;
   30579: out<=0;
   30580: out<=1;
   30581: out<=1;
   30582: out<=1;
   30583: out<=1;
   30584: out<=1;
   30585: out<=1;
   30586: out<=0;
   30587: out<=0;
   30588: out<=0;
   30589: out<=1;
   30590: out<=0;
   30591: out<=1;
   30592: out<=1;
   30593: out<=0;
   30594: out<=0;
   30595: out<=1;
   30596: out<=0;
   30597: out<=0;
   30598: out<=0;
   30599: out<=0;
   30600: out<=0;
   30601: out<=0;
   30602: out<=1;
   30603: out<=1;
   30604: out<=1;
   30605: out<=0;
   30606: out<=1;
   30607: out<=0;
   30608: out<=0;
   30609: out<=1;
   30610: out<=1;
   30611: out<=0;
   30612: out<=1;
   30613: out<=1;
   30614: out<=1;
   30615: out<=1;
   30616: out<=1;
   30617: out<=1;
   30618: out<=0;
   30619: out<=0;
   30620: out<=0;
   30621: out<=1;
   30622: out<=0;
   30623: out<=1;
   30624: out<=0;
   30625: out<=1;
   30626: out<=1;
   30627: out<=0;
   30628: out<=1;
   30629: out<=1;
   30630: out<=1;
   30631: out<=1;
   30632: out<=1;
   30633: out<=1;
   30634: out<=0;
   30635: out<=0;
   30636: out<=0;
   30637: out<=1;
   30638: out<=0;
   30639: out<=1;
   30640: out<=1;
   30641: out<=0;
   30642: out<=0;
   30643: out<=1;
   30644: out<=0;
   30645: out<=0;
   30646: out<=0;
   30647: out<=0;
   30648: out<=0;
   30649: out<=0;
   30650: out<=1;
   30651: out<=1;
   30652: out<=1;
   30653: out<=0;
   30654: out<=1;
   30655: out<=0;
   30656: out<=0;
   30657: out<=1;
   30658: out<=1;
   30659: out<=0;
   30660: out<=1;
   30661: out<=1;
   30662: out<=1;
   30663: out<=1;
   30664: out<=1;
   30665: out<=1;
   30666: out<=0;
   30667: out<=0;
   30668: out<=0;
   30669: out<=1;
   30670: out<=0;
   30671: out<=1;
   30672: out<=0;
   30673: out<=1;
   30674: out<=1;
   30675: out<=0;
   30676: out<=1;
   30677: out<=1;
   30678: out<=1;
   30679: out<=1;
   30680: out<=1;
   30681: out<=1;
   30682: out<=0;
   30683: out<=0;
   30684: out<=0;
   30685: out<=1;
   30686: out<=0;
   30687: out<=1;
   30688: out<=0;
   30689: out<=1;
   30690: out<=1;
   30691: out<=0;
   30692: out<=1;
   30693: out<=1;
   30694: out<=1;
   30695: out<=1;
   30696: out<=1;
   30697: out<=1;
   30698: out<=0;
   30699: out<=0;
   30700: out<=0;
   30701: out<=1;
   30702: out<=0;
   30703: out<=1;
   30704: out<=0;
   30705: out<=1;
   30706: out<=1;
   30707: out<=0;
   30708: out<=1;
   30709: out<=1;
   30710: out<=1;
   30711: out<=1;
   30712: out<=1;
   30713: out<=1;
   30714: out<=0;
   30715: out<=0;
   30716: out<=0;
   30717: out<=1;
   30718: out<=0;
   30719: out<=1;
   30720: out<=0;
   30721: out<=1;
   30722: out<=1;
   30723: out<=0;
   30724: out<=1;
   30725: out<=1;
   30726: out<=1;
   30727: out<=1;
   30728: out<=0;
   30729: out<=0;
   30730: out<=1;
   30731: out<=1;
   30732: out<=1;
   30733: out<=0;
   30734: out<=1;
   30735: out<=0;
   30736: out<=0;
   30737: out<=1;
   30738: out<=1;
   30739: out<=0;
   30740: out<=1;
   30741: out<=1;
   30742: out<=1;
   30743: out<=1;
   30744: out<=0;
   30745: out<=0;
   30746: out<=1;
   30747: out<=1;
   30748: out<=1;
   30749: out<=0;
   30750: out<=1;
   30751: out<=0;
   30752: out<=0;
   30753: out<=1;
   30754: out<=1;
   30755: out<=0;
   30756: out<=1;
   30757: out<=1;
   30758: out<=1;
   30759: out<=1;
   30760: out<=0;
   30761: out<=0;
   30762: out<=1;
   30763: out<=1;
   30764: out<=1;
   30765: out<=0;
   30766: out<=1;
   30767: out<=0;
   30768: out<=0;
   30769: out<=1;
   30770: out<=1;
   30771: out<=0;
   30772: out<=1;
   30773: out<=1;
   30774: out<=1;
   30775: out<=1;
   30776: out<=0;
   30777: out<=0;
   30778: out<=1;
   30779: out<=1;
   30780: out<=1;
   30781: out<=0;
   30782: out<=1;
   30783: out<=0;
   30784: out<=1;
   30785: out<=0;
   30786: out<=0;
   30787: out<=1;
   30788: out<=0;
   30789: out<=0;
   30790: out<=0;
   30791: out<=0;
   30792: out<=1;
   30793: out<=1;
   30794: out<=0;
   30795: out<=0;
   30796: out<=0;
   30797: out<=1;
   30798: out<=0;
   30799: out<=1;
   30800: out<=0;
   30801: out<=1;
   30802: out<=1;
   30803: out<=0;
   30804: out<=1;
   30805: out<=1;
   30806: out<=1;
   30807: out<=1;
   30808: out<=0;
   30809: out<=0;
   30810: out<=1;
   30811: out<=1;
   30812: out<=1;
   30813: out<=0;
   30814: out<=1;
   30815: out<=0;
   30816: out<=0;
   30817: out<=1;
   30818: out<=1;
   30819: out<=0;
   30820: out<=1;
   30821: out<=1;
   30822: out<=1;
   30823: out<=1;
   30824: out<=0;
   30825: out<=0;
   30826: out<=1;
   30827: out<=1;
   30828: out<=1;
   30829: out<=0;
   30830: out<=1;
   30831: out<=0;
   30832: out<=1;
   30833: out<=0;
   30834: out<=0;
   30835: out<=1;
   30836: out<=0;
   30837: out<=0;
   30838: out<=0;
   30839: out<=0;
   30840: out<=1;
   30841: out<=1;
   30842: out<=0;
   30843: out<=0;
   30844: out<=0;
   30845: out<=1;
   30846: out<=0;
   30847: out<=1;
   30848: out<=1;
   30849: out<=0;
   30850: out<=0;
   30851: out<=1;
   30852: out<=0;
   30853: out<=0;
   30854: out<=0;
   30855: out<=0;
   30856: out<=1;
   30857: out<=1;
   30858: out<=0;
   30859: out<=0;
   30860: out<=0;
   30861: out<=1;
   30862: out<=0;
   30863: out<=1;
   30864: out<=0;
   30865: out<=1;
   30866: out<=1;
   30867: out<=0;
   30868: out<=1;
   30869: out<=1;
   30870: out<=1;
   30871: out<=1;
   30872: out<=0;
   30873: out<=0;
   30874: out<=1;
   30875: out<=1;
   30876: out<=1;
   30877: out<=0;
   30878: out<=1;
   30879: out<=0;
   30880: out<=1;
   30881: out<=0;
   30882: out<=0;
   30883: out<=1;
   30884: out<=0;
   30885: out<=0;
   30886: out<=0;
   30887: out<=0;
   30888: out<=1;
   30889: out<=1;
   30890: out<=0;
   30891: out<=0;
   30892: out<=0;
   30893: out<=1;
   30894: out<=0;
   30895: out<=1;
   30896: out<=0;
   30897: out<=1;
   30898: out<=1;
   30899: out<=0;
   30900: out<=1;
   30901: out<=1;
   30902: out<=1;
   30903: out<=1;
   30904: out<=0;
   30905: out<=0;
   30906: out<=1;
   30907: out<=1;
   30908: out<=1;
   30909: out<=0;
   30910: out<=1;
   30911: out<=0;
   30912: out<=0;
   30913: out<=1;
   30914: out<=1;
   30915: out<=0;
   30916: out<=1;
   30917: out<=1;
   30918: out<=1;
   30919: out<=1;
   30920: out<=0;
   30921: out<=0;
   30922: out<=1;
   30923: out<=1;
   30924: out<=1;
   30925: out<=0;
   30926: out<=1;
   30927: out<=0;
   30928: out<=0;
   30929: out<=1;
   30930: out<=1;
   30931: out<=0;
   30932: out<=1;
   30933: out<=1;
   30934: out<=1;
   30935: out<=1;
   30936: out<=0;
   30937: out<=0;
   30938: out<=1;
   30939: out<=1;
   30940: out<=1;
   30941: out<=0;
   30942: out<=1;
   30943: out<=0;
   30944: out<=1;
   30945: out<=0;
   30946: out<=0;
   30947: out<=1;
   30948: out<=0;
   30949: out<=0;
   30950: out<=0;
   30951: out<=0;
   30952: out<=1;
   30953: out<=1;
   30954: out<=0;
   30955: out<=0;
   30956: out<=0;
   30957: out<=1;
   30958: out<=0;
   30959: out<=1;
   30960: out<=1;
   30961: out<=0;
   30962: out<=0;
   30963: out<=1;
   30964: out<=0;
   30965: out<=0;
   30966: out<=0;
   30967: out<=0;
   30968: out<=1;
   30969: out<=1;
   30970: out<=0;
   30971: out<=0;
   30972: out<=0;
   30973: out<=1;
   30974: out<=0;
   30975: out<=1;
   30976: out<=1;
   30977: out<=1;
   30978: out<=1;
   30979: out<=1;
   30980: out<=1;
   30981: out<=0;
   30982: out<=0;
   30983: out<=1;
   30984: out<=0;
   30985: out<=1;
   30986: out<=0;
   30987: out<=1;
   30988: out<=0;
   30989: out<=0;
   30990: out<=1;
   30991: out<=1;
   30992: out<=0;
   30993: out<=0;
   30994: out<=0;
   30995: out<=0;
   30996: out<=0;
   30997: out<=1;
   30998: out<=1;
   30999: out<=0;
   31000: out<=1;
   31001: out<=0;
   31002: out<=1;
   31003: out<=0;
   31004: out<=1;
   31005: out<=1;
   31006: out<=0;
   31007: out<=0;
   31008: out<=0;
   31009: out<=0;
   31010: out<=0;
   31011: out<=0;
   31012: out<=0;
   31013: out<=1;
   31014: out<=1;
   31015: out<=0;
   31016: out<=1;
   31017: out<=0;
   31018: out<=1;
   31019: out<=0;
   31020: out<=1;
   31021: out<=1;
   31022: out<=0;
   31023: out<=0;
   31024: out<=1;
   31025: out<=1;
   31026: out<=1;
   31027: out<=1;
   31028: out<=1;
   31029: out<=0;
   31030: out<=0;
   31031: out<=1;
   31032: out<=0;
   31033: out<=1;
   31034: out<=0;
   31035: out<=1;
   31036: out<=0;
   31037: out<=0;
   31038: out<=1;
   31039: out<=1;
   31040: out<=0;
   31041: out<=0;
   31042: out<=0;
   31043: out<=0;
   31044: out<=0;
   31045: out<=1;
   31046: out<=1;
   31047: out<=0;
   31048: out<=1;
   31049: out<=0;
   31050: out<=1;
   31051: out<=0;
   31052: out<=1;
   31053: out<=1;
   31054: out<=0;
   31055: out<=0;
   31056: out<=0;
   31057: out<=0;
   31058: out<=0;
   31059: out<=0;
   31060: out<=0;
   31061: out<=1;
   31062: out<=1;
   31063: out<=0;
   31064: out<=1;
   31065: out<=0;
   31066: out<=1;
   31067: out<=0;
   31068: out<=1;
   31069: out<=1;
   31070: out<=0;
   31071: out<=0;
   31072: out<=0;
   31073: out<=0;
   31074: out<=0;
   31075: out<=0;
   31076: out<=0;
   31077: out<=1;
   31078: out<=1;
   31079: out<=0;
   31080: out<=1;
   31081: out<=0;
   31082: out<=1;
   31083: out<=0;
   31084: out<=1;
   31085: out<=1;
   31086: out<=0;
   31087: out<=0;
   31088: out<=0;
   31089: out<=0;
   31090: out<=0;
   31091: out<=0;
   31092: out<=0;
   31093: out<=1;
   31094: out<=1;
   31095: out<=0;
   31096: out<=1;
   31097: out<=0;
   31098: out<=1;
   31099: out<=0;
   31100: out<=1;
   31101: out<=1;
   31102: out<=0;
   31103: out<=0;
   31104: out<=0;
   31105: out<=0;
   31106: out<=0;
   31107: out<=0;
   31108: out<=0;
   31109: out<=1;
   31110: out<=1;
   31111: out<=0;
   31112: out<=1;
   31113: out<=0;
   31114: out<=1;
   31115: out<=0;
   31116: out<=1;
   31117: out<=1;
   31118: out<=0;
   31119: out<=0;
   31120: out<=0;
   31121: out<=0;
   31122: out<=0;
   31123: out<=0;
   31124: out<=0;
   31125: out<=1;
   31126: out<=1;
   31127: out<=0;
   31128: out<=1;
   31129: out<=0;
   31130: out<=1;
   31131: out<=0;
   31132: out<=1;
   31133: out<=1;
   31134: out<=0;
   31135: out<=0;
   31136: out<=1;
   31137: out<=1;
   31138: out<=1;
   31139: out<=1;
   31140: out<=1;
   31141: out<=0;
   31142: out<=0;
   31143: out<=1;
   31144: out<=0;
   31145: out<=1;
   31146: out<=0;
   31147: out<=1;
   31148: out<=0;
   31149: out<=0;
   31150: out<=1;
   31151: out<=1;
   31152: out<=1;
   31153: out<=1;
   31154: out<=1;
   31155: out<=1;
   31156: out<=1;
   31157: out<=0;
   31158: out<=0;
   31159: out<=1;
   31160: out<=0;
   31161: out<=1;
   31162: out<=0;
   31163: out<=1;
   31164: out<=0;
   31165: out<=0;
   31166: out<=1;
   31167: out<=1;
   31168: out<=1;
   31169: out<=1;
   31170: out<=1;
   31171: out<=1;
   31172: out<=1;
   31173: out<=0;
   31174: out<=0;
   31175: out<=1;
   31176: out<=0;
   31177: out<=1;
   31178: out<=0;
   31179: out<=1;
   31180: out<=0;
   31181: out<=0;
   31182: out<=1;
   31183: out<=1;
   31184: out<=0;
   31185: out<=0;
   31186: out<=0;
   31187: out<=0;
   31188: out<=0;
   31189: out<=1;
   31190: out<=1;
   31191: out<=0;
   31192: out<=1;
   31193: out<=0;
   31194: out<=1;
   31195: out<=0;
   31196: out<=1;
   31197: out<=1;
   31198: out<=0;
   31199: out<=0;
   31200: out<=1;
   31201: out<=1;
   31202: out<=1;
   31203: out<=1;
   31204: out<=1;
   31205: out<=0;
   31206: out<=0;
   31207: out<=1;
   31208: out<=0;
   31209: out<=1;
   31210: out<=0;
   31211: out<=1;
   31212: out<=0;
   31213: out<=0;
   31214: out<=1;
   31215: out<=1;
   31216: out<=0;
   31217: out<=0;
   31218: out<=0;
   31219: out<=0;
   31220: out<=0;
   31221: out<=1;
   31222: out<=1;
   31223: out<=0;
   31224: out<=1;
   31225: out<=0;
   31226: out<=1;
   31227: out<=0;
   31228: out<=1;
   31229: out<=1;
   31230: out<=0;
   31231: out<=0;
   31232: out<=0;
   31233: out<=0;
   31234: out<=1;
   31235: out<=1;
   31236: out<=0;
   31237: out<=1;
   31238: out<=0;
   31239: out<=1;
   31240: out<=0;
   31241: out<=1;
   31242: out<=1;
   31243: out<=0;
   31244: out<=0;
   31245: out<=0;
   31246: out<=0;
   31247: out<=0;
   31248: out<=1;
   31249: out<=1;
   31250: out<=0;
   31251: out<=0;
   31252: out<=1;
   31253: out<=0;
   31254: out<=1;
   31255: out<=0;
   31256: out<=1;
   31257: out<=0;
   31258: out<=0;
   31259: out<=1;
   31260: out<=1;
   31261: out<=1;
   31262: out<=1;
   31263: out<=1;
   31264: out<=0;
   31265: out<=0;
   31266: out<=1;
   31267: out<=1;
   31268: out<=0;
   31269: out<=1;
   31270: out<=0;
   31271: out<=1;
   31272: out<=0;
   31273: out<=1;
   31274: out<=1;
   31275: out<=0;
   31276: out<=0;
   31277: out<=0;
   31278: out<=0;
   31279: out<=0;
   31280: out<=1;
   31281: out<=1;
   31282: out<=0;
   31283: out<=0;
   31284: out<=1;
   31285: out<=0;
   31286: out<=1;
   31287: out<=0;
   31288: out<=1;
   31289: out<=0;
   31290: out<=0;
   31291: out<=1;
   31292: out<=1;
   31293: out<=1;
   31294: out<=1;
   31295: out<=1;
   31296: out<=1;
   31297: out<=1;
   31298: out<=0;
   31299: out<=0;
   31300: out<=1;
   31301: out<=0;
   31302: out<=1;
   31303: out<=0;
   31304: out<=1;
   31305: out<=0;
   31306: out<=0;
   31307: out<=1;
   31308: out<=1;
   31309: out<=1;
   31310: out<=1;
   31311: out<=1;
   31312: out<=1;
   31313: out<=1;
   31314: out<=0;
   31315: out<=0;
   31316: out<=1;
   31317: out<=0;
   31318: out<=1;
   31319: out<=0;
   31320: out<=1;
   31321: out<=0;
   31322: out<=0;
   31323: out<=1;
   31324: out<=1;
   31325: out<=1;
   31326: out<=1;
   31327: out<=1;
   31328: out<=0;
   31329: out<=0;
   31330: out<=1;
   31331: out<=1;
   31332: out<=0;
   31333: out<=1;
   31334: out<=0;
   31335: out<=1;
   31336: out<=0;
   31337: out<=1;
   31338: out<=1;
   31339: out<=0;
   31340: out<=0;
   31341: out<=0;
   31342: out<=0;
   31343: out<=0;
   31344: out<=0;
   31345: out<=0;
   31346: out<=1;
   31347: out<=1;
   31348: out<=0;
   31349: out<=1;
   31350: out<=0;
   31351: out<=1;
   31352: out<=0;
   31353: out<=1;
   31354: out<=1;
   31355: out<=0;
   31356: out<=0;
   31357: out<=0;
   31358: out<=0;
   31359: out<=0;
   31360: out<=1;
   31361: out<=1;
   31362: out<=0;
   31363: out<=0;
   31364: out<=1;
   31365: out<=0;
   31366: out<=1;
   31367: out<=0;
   31368: out<=1;
   31369: out<=0;
   31370: out<=0;
   31371: out<=1;
   31372: out<=1;
   31373: out<=1;
   31374: out<=1;
   31375: out<=1;
   31376: out<=1;
   31377: out<=1;
   31378: out<=0;
   31379: out<=0;
   31380: out<=1;
   31381: out<=0;
   31382: out<=1;
   31383: out<=0;
   31384: out<=1;
   31385: out<=0;
   31386: out<=0;
   31387: out<=1;
   31388: out<=1;
   31389: out<=1;
   31390: out<=1;
   31391: out<=1;
   31392: out<=1;
   31393: out<=1;
   31394: out<=0;
   31395: out<=0;
   31396: out<=1;
   31397: out<=0;
   31398: out<=1;
   31399: out<=0;
   31400: out<=1;
   31401: out<=0;
   31402: out<=0;
   31403: out<=1;
   31404: out<=1;
   31405: out<=1;
   31406: out<=1;
   31407: out<=1;
   31408: out<=1;
   31409: out<=1;
   31410: out<=0;
   31411: out<=0;
   31412: out<=1;
   31413: out<=0;
   31414: out<=1;
   31415: out<=0;
   31416: out<=1;
   31417: out<=0;
   31418: out<=0;
   31419: out<=1;
   31420: out<=1;
   31421: out<=1;
   31422: out<=1;
   31423: out<=1;
   31424: out<=0;
   31425: out<=0;
   31426: out<=1;
   31427: out<=1;
   31428: out<=0;
   31429: out<=1;
   31430: out<=0;
   31431: out<=1;
   31432: out<=0;
   31433: out<=1;
   31434: out<=1;
   31435: out<=0;
   31436: out<=0;
   31437: out<=0;
   31438: out<=0;
   31439: out<=0;
   31440: out<=1;
   31441: out<=1;
   31442: out<=0;
   31443: out<=0;
   31444: out<=1;
   31445: out<=0;
   31446: out<=1;
   31447: out<=0;
   31448: out<=1;
   31449: out<=0;
   31450: out<=0;
   31451: out<=1;
   31452: out<=1;
   31453: out<=1;
   31454: out<=1;
   31455: out<=1;
   31456: out<=1;
   31457: out<=1;
   31458: out<=0;
   31459: out<=0;
   31460: out<=1;
   31461: out<=0;
   31462: out<=1;
   31463: out<=0;
   31464: out<=1;
   31465: out<=0;
   31466: out<=0;
   31467: out<=1;
   31468: out<=1;
   31469: out<=1;
   31470: out<=1;
   31471: out<=1;
   31472: out<=0;
   31473: out<=0;
   31474: out<=1;
   31475: out<=1;
   31476: out<=0;
   31477: out<=1;
   31478: out<=0;
   31479: out<=1;
   31480: out<=0;
   31481: out<=1;
   31482: out<=1;
   31483: out<=0;
   31484: out<=0;
   31485: out<=0;
   31486: out<=0;
   31487: out<=0;
   31488: out<=1;
   31489: out<=0;
   31490: out<=1;
   31491: out<=0;
   31492: out<=0;
   31493: out<=0;
   31494: out<=1;
   31495: out<=1;
   31496: out<=0;
   31497: out<=0;
   31498: out<=0;
   31499: out<=0;
   31500: out<=1;
   31501: out<=0;
   31502: out<=0;
   31503: out<=1;
   31504: out<=1;
   31505: out<=0;
   31506: out<=1;
   31507: out<=0;
   31508: out<=0;
   31509: out<=0;
   31510: out<=1;
   31511: out<=1;
   31512: out<=0;
   31513: out<=0;
   31514: out<=0;
   31515: out<=0;
   31516: out<=1;
   31517: out<=0;
   31518: out<=0;
   31519: out<=1;
   31520: out<=0;
   31521: out<=1;
   31522: out<=0;
   31523: out<=1;
   31524: out<=1;
   31525: out<=1;
   31526: out<=0;
   31527: out<=0;
   31528: out<=1;
   31529: out<=1;
   31530: out<=1;
   31531: out<=1;
   31532: out<=0;
   31533: out<=1;
   31534: out<=1;
   31535: out<=0;
   31536: out<=0;
   31537: out<=1;
   31538: out<=0;
   31539: out<=1;
   31540: out<=1;
   31541: out<=1;
   31542: out<=0;
   31543: out<=0;
   31544: out<=1;
   31545: out<=1;
   31546: out<=1;
   31547: out<=1;
   31548: out<=0;
   31549: out<=1;
   31550: out<=1;
   31551: out<=0;
   31552: out<=0;
   31553: out<=1;
   31554: out<=0;
   31555: out<=1;
   31556: out<=1;
   31557: out<=1;
   31558: out<=0;
   31559: out<=0;
   31560: out<=1;
   31561: out<=1;
   31562: out<=1;
   31563: out<=1;
   31564: out<=0;
   31565: out<=1;
   31566: out<=1;
   31567: out<=0;
   31568: out<=1;
   31569: out<=0;
   31570: out<=1;
   31571: out<=0;
   31572: out<=0;
   31573: out<=0;
   31574: out<=1;
   31575: out<=1;
   31576: out<=0;
   31577: out<=0;
   31578: out<=0;
   31579: out<=0;
   31580: out<=1;
   31581: out<=0;
   31582: out<=0;
   31583: out<=1;
   31584: out<=0;
   31585: out<=1;
   31586: out<=0;
   31587: out<=1;
   31588: out<=1;
   31589: out<=1;
   31590: out<=0;
   31591: out<=0;
   31592: out<=1;
   31593: out<=1;
   31594: out<=1;
   31595: out<=1;
   31596: out<=0;
   31597: out<=1;
   31598: out<=1;
   31599: out<=0;
   31600: out<=1;
   31601: out<=0;
   31602: out<=1;
   31603: out<=0;
   31604: out<=0;
   31605: out<=0;
   31606: out<=1;
   31607: out<=1;
   31608: out<=0;
   31609: out<=0;
   31610: out<=0;
   31611: out<=0;
   31612: out<=1;
   31613: out<=0;
   31614: out<=0;
   31615: out<=1;
   31616: out<=0;
   31617: out<=1;
   31618: out<=0;
   31619: out<=1;
   31620: out<=1;
   31621: out<=1;
   31622: out<=0;
   31623: out<=0;
   31624: out<=1;
   31625: out<=1;
   31626: out<=1;
   31627: out<=1;
   31628: out<=0;
   31629: out<=1;
   31630: out<=1;
   31631: out<=0;
   31632: out<=1;
   31633: out<=0;
   31634: out<=1;
   31635: out<=0;
   31636: out<=0;
   31637: out<=0;
   31638: out<=1;
   31639: out<=1;
   31640: out<=0;
   31641: out<=0;
   31642: out<=0;
   31643: out<=0;
   31644: out<=1;
   31645: out<=0;
   31646: out<=0;
   31647: out<=1;
   31648: out<=1;
   31649: out<=0;
   31650: out<=1;
   31651: out<=0;
   31652: out<=0;
   31653: out<=0;
   31654: out<=1;
   31655: out<=1;
   31656: out<=0;
   31657: out<=0;
   31658: out<=0;
   31659: out<=0;
   31660: out<=1;
   31661: out<=0;
   31662: out<=0;
   31663: out<=1;
   31664: out<=0;
   31665: out<=1;
   31666: out<=0;
   31667: out<=1;
   31668: out<=1;
   31669: out<=1;
   31670: out<=0;
   31671: out<=0;
   31672: out<=1;
   31673: out<=1;
   31674: out<=1;
   31675: out<=1;
   31676: out<=0;
   31677: out<=1;
   31678: out<=1;
   31679: out<=0;
   31680: out<=1;
   31681: out<=0;
   31682: out<=1;
   31683: out<=0;
   31684: out<=0;
   31685: out<=0;
   31686: out<=1;
   31687: out<=1;
   31688: out<=0;
   31689: out<=0;
   31690: out<=0;
   31691: out<=0;
   31692: out<=1;
   31693: out<=0;
   31694: out<=0;
   31695: out<=1;
   31696: out<=1;
   31697: out<=0;
   31698: out<=1;
   31699: out<=0;
   31700: out<=0;
   31701: out<=0;
   31702: out<=1;
   31703: out<=1;
   31704: out<=0;
   31705: out<=0;
   31706: out<=0;
   31707: out<=0;
   31708: out<=1;
   31709: out<=0;
   31710: out<=0;
   31711: out<=1;
   31712: out<=1;
   31713: out<=0;
   31714: out<=1;
   31715: out<=0;
   31716: out<=0;
   31717: out<=0;
   31718: out<=1;
   31719: out<=1;
   31720: out<=0;
   31721: out<=0;
   31722: out<=0;
   31723: out<=0;
   31724: out<=1;
   31725: out<=0;
   31726: out<=0;
   31727: out<=1;
   31728: out<=1;
   31729: out<=0;
   31730: out<=1;
   31731: out<=0;
   31732: out<=0;
   31733: out<=0;
   31734: out<=1;
   31735: out<=1;
   31736: out<=0;
   31737: out<=0;
   31738: out<=0;
   31739: out<=0;
   31740: out<=1;
   31741: out<=0;
   31742: out<=0;
   31743: out<=1;
   31744: out<=0;
   31745: out<=0;
   31746: out<=0;
   31747: out<=0;
   31748: out<=1;
   31749: out<=0;
   31750: out<=0;
   31751: out<=1;
   31752: out<=0;
   31753: out<=1;
   31754: out<=0;
   31755: out<=1;
   31756: out<=1;
   31757: out<=1;
   31758: out<=0;
   31759: out<=0;
   31760: out<=0;
   31761: out<=0;
   31762: out<=0;
   31763: out<=0;
   31764: out<=1;
   31765: out<=0;
   31766: out<=0;
   31767: out<=1;
   31768: out<=0;
   31769: out<=1;
   31770: out<=0;
   31771: out<=1;
   31772: out<=1;
   31773: out<=1;
   31774: out<=0;
   31775: out<=0;
   31776: out<=0;
   31777: out<=0;
   31778: out<=0;
   31779: out<=0;
   31780: out<=1;
   31781: out<=0;
   31782: out<=0;
   31783: out<=1;
   31784: out<=0;
   31785: out<=1;
   31786: out<=0;
   31787: out<=1;
   31788: out<=1;
   31789: out<=1;
   31790: out<=0;
   31791: out<=0;
   31792: out<=0;
   31793: out<=0;
   31794: out<=0;
   31795: out<=0;
   31796: out<=1;
   31797: out<=0;
   31798: out<=0;
   31799: out<=1;
   31800: out<=0;
   31801: out<=1;
   31802: out<=0;
   31803: out<=1;
   31804: out<=1;
   31805: out<=1;
   31806: out<=0;
   31807: out<=0;
   31808: out<=1;
   31809: out<=1;
   31810: out<=1;
   31811: out<=1;
   31812: out<=0;
   31813: out<=1;
   31814: out<=1;
   31815: out<=0;
   31816: out<=1;
   31817: out<=0;
   31818: out<=1;
   31819: out<=0;
   31820: out<=0;
   31821: out<=0;
   31822: out<=1;
   31823: out<=1;
   31824: out<=0;
   31825: out<=0;
   31826: out<=0;
   31827: out<=0;
   31828: out<=1;
   31829: out<=0;
   31830: out<=0;
   31831: out<=1;
   31832: out<=0;
   31833: out<=1;
   31834: out<=0;
   31835: out<=1;
   31836: out<=1;
   31837: out<=1;
   31838: out<=0;
   31839: out<=0;
   31840: out<=0;
   31841: out<=0;
   31842: out<=0;
   31843: out<=0;
   31844: out<=1;
   31845: out<=0;
   31846: out<=0;
   31847: out<=1;
   31848: out<=0;
   31849: out<=1;
   31850: out<=0;
   31851: out<=1;
   31852: out<=1;
   31853: out<=1;
   31854: out<=0;
   31855: out<=0;
   31856: out<=1;
   31857: out<=1;
   31858: out<=1;
   31859: out<=1;
   31860: out<=0;
   31861: out<=1;
   31862: out<=1;
   31863: out<=0;
   31864: out<=1;
   31865: out<=0;
   31866: out<=1;
   31867: out<=0;
   31868: out<=0;
   31869: out<=0;
   31870: out<=1;
   31871: out<=1;
   31872: out<=1;
   31873: out<=1;
   31874: out<=1;
   31875: out<=1;
   31876: out<=0;
   31877: out<=1;
   31878: out<=1;
   31879: out<=0;
   31880: out<=1;
   31881: out<=0;
   31882: out<=1;
   31883: out<=0;
   31884: out<=0;
   31885: out<=0;
   31886: out<=1;
   31887: out<=1;
   31888: out<=0;
   31889: out<=0;
   31890: out<=0;
   31891: out<=0;
   31892: out<=1;
   31893: out<=0;
   31894: out<=0;
   31895: out<=1;
   31896: out<=0;
   31897: out<=1;
   31898: out<=0;
   31899: out<=1;
   31900: out<=1;
   31901: out<=1;
   31902: out<=0;
   31903: out<=0;
   31904: out<=1;
   31905: out<=1;
   31906: out<=1;
   31907: out<=1;
   31908: out<=0;
   31909: out<=1;
   31910: out<=1;
   31911: out<=0;
   31912: out<=1;
   31913: out<=0;
   31914: out<=1;
   31915: out<=0;
   31916: out<=0;
   31917: out<=0;
   31918: out<=1;
   31919: out<=1;
   31920: out<=0;
   31921: out<=0;
   31922: out<=0;
   31923: out<=0;
   31924: out<=1;
   31925: out<=0;
   31926: out<=0;
   31927: out<=1;
   31928: out<=0;
   31929: out<=1;
   31930: out<=0;
   31931: out<=1;
   31932: out<=1;
   31933: out<=1;
   31934: out<=0;
   31935: out<=0;
   31936: out<=0;
   31937: out<=0;
   31938: out<=0;
   31939: out<=0;
   31940: out<=1;
   31941: out<=0;
   31942: out<=0;
   31943: out<=1;
   31944: out<=0;
   31945: out<=1;
   31946: out<=0;
   31947: out<=1;
   31948: out<=1;
   31949: out<=1;
   31950: out<=0;
   31951: out<=0;
   31952: out<=0;
   31953: out<=0;
   31954: out<=0;
   31955: out<=0;
   31956: out<=1;
   31957: out<=0;
   31958: out<=0;
   31959: out<=1;
   31960: out<=0;
   31961: out<=1;
   31962: out<=0;
   31963: out<=1;
   31964: out<=1;
   31965: out<=1;
   31966: out<=0;
   31967: out<=0;
   31968: out<=1;
   31969: out<=1;
   31970: out<=1;
   31971: out<=1;
   31972: out<=0;
   31973: out<=1;
   31974: out<=1;
   31975: out<=0;
   31976: out<=1;
   31977: out<=0;
   31978: out<=1;
   31979: out<=0;
   31980: out<=0;
   31981: out<=0;
   31982: out<=1;
   31983: out<=1;
   31984: out<=1;
   31985: out<=1;
   31986: out<=1;
   31987: out<=1;
   31988: out<=0;
   31989: out<=1;
   31990: out<=1;
   31991: out<=0;
   31992: out<=1;
   31993: out<=0;
   31994: out<=1;
   31995: out<=0;
   31996: out<=0;
   31997: out<=0;
   31998: out<=1;
   31999: out<=1;
   32000: out<=0;
   32001: out<=1;
   32002: out<=1;
   32003: out<=0;
   32004: out<=0;
   32005: out<=0;
   32006: out<=0;
   32007: out<=0;
   32008: out<=1;
   32009: out<=1;
   32010: out<=0;
   32011: out<=0;
   32012: out<=1;
   32013: out<=0;
   32014: out<=1;
   32015: out<=0;
   32016: out<=1;
   32017: out<=0;
   32018: out<=0;
   32019: out<=1;
   32020: out<=1;
   32021: out<=1;
   32022: out<=1;
   32023: out<=1;
   32024: out<=0;
   32025: out<=0;
   32026: out<=1;
   32027: out<=1;
   32028: out<=0;
   32029: out<=1;
   32030: out<=0;
   32031: out<=1;
   32032: out<=1;
   32033: out<=0;
   32034: out<=0;
   32035: out<=1;
   32036: out<=1;
   32037: out<=1;
   32038: out<=1;
   32039: out<=1;
   32040: out<=0;
   32041: out<=0;
   32042: out<=1;
   32043: out<=1;
   32044: out<=0;
   32045: out<=1;
   32046: out<=0;
   32047: out<=1;
   32048: out<=0;
   32049: out<=1;
   32050: out<=1;
   32051: out<=0;
   32052: out<=0;
   32053: out<=0;
   32054: out<=0;
   32055: out<=0;
   32056: out<=1;
   32057: out<=1;
   32058: out<=0;
   32059: out<=0;
   32060: out<=1;
   32061: out<=0;
   32062: out<=1;
   32063: out<=0;
   32064: out<=1;
   32065: out<=0;
   32066: out<=0;
   32067: out<=1;
   32068: out<=1;
   32069: out<=1;
   32070: out<=1;
   32071: out<=1;
   32072: out<=0;
   32073: out<=0;
   32074: out<=1;
   32075: out<=1;
   32076: out<=0;
   32077: out<=1;
   32078: out<=0;
   32079: out<=1;
   32080: out<=1;
   32081: out<=0;
   32082: out<=0;
   32083: out<=1;
   32084: out<=1;
   32085: out<=1;
   32086: out<=1;
   32087: out<=1;
   32088: out<=0;
   32089: out<=0;
   32090: out<=1;
   32091: out<=1;
   32092: out<=0;
   32093: out<=1;
   32094: out<=0;
   32095: out<=1;
   32096: out<=1;
   32097: out<=0;
   32098: out<=0;
   32099: out<=1;
   32100: out<=1;
   32101: out<=1;
   32102: out<=1;
   32103: out<=1;
   32104: out<=0;
   32105: out<=0;
   32106: out<=1;
   32107: out<=1;
   32108: out<=0;
   32109: out<=1;
   32110: out<=0;
   32111: out<=1;
   32112: out<=1;
   32113: out<=0;
   32114: out<=0;
   32115: out<=1;
   32116: out<=1;
   32117: out<=1;
   32118: out<=1;
   32119: out<=1;
   32120: out<=0;
   32121: out<=0;
   32122: out<=1;
   32123: out<=1;
   32124: out<=0;
   32125: out<=1;
   32126: out<=0;
   32127: out<=1;
   32128: out<=1;
   32129: out<=0;
   32130: out<=0;
   32131: out<=1;
   32132: out<=1;
   32133: out<=1;
   32134: out<=1;
   32135: out<=1;
   32136: out<=0;
   32137: out<=0;
   32138: out<=1;
   32139: out<=1;
   32140: out<=0;
   32141: out<=1;
   32142: out<=0;
   32143: out<=1;
   32144: out<=1;
   32145: out<=0;
   32146: out<=0;
   32147: out<=1;
   32148: out<=1;
   32149: out<=1;
   32150: out<=1;
   32151: out<=1;
   32152: out<=0;
   32153: out<=0;
   32154: out<=1;
   32155: out<=1;
   32156: out<=0;
   32157: out<=1;
   32158: out<=0;
   32159: out<=1;
   32160: out<=0;
   32161: out<=1;
   32162: out<=1;
   32163: out<=0;
   32164: out<=0;
   32165: out<=0;
   32166: out<=0;
   32167: out<=0;
   32168: out<=1;
   32169: out<=1;
   32170: out<=0;
   32171: out<=0;
   32172: out<=1;
   32173: out<=0;
   32174: out<=1;
   32175: out<=0;
   32176: out<=0;
   32177: out<=1;
   32178: out<=1;
   32179: out<=0;
   32180: out<=0;
   32181: out<=0;
   32182: out<=0;
   32183: out<=0;
   32184: out<=1;
   32185: out<=1;
   32186: out<=0;
   32187: out<=0;
   32188: out<=1;
   32189: out<=0;
   32190: out<=1;
   32191: out<=0;
   32192: out<=0;
   32193: out<=1;
   32194: out<=1;
   32195: out<=0;
   32196: out<=0;
   32197: out<=0;
   32198: out<=0;
   32199: out<=0;
   32200: out<=1;
   32201: out<=1;
   32202: out<=0;
   32203: out<=0;
   32204: out<=1;
   32205: out<=0;
   32206: out<=1;
   32207: out<=0;
   32208: out<=1;
   32209: out<=0;
   32210: out<=0;
   32211: out<=1;
   32212: out<=1;
   32213: out<=1;
   32214: out<=1;
   32215: out<=1;
   32216: out<=0;
   32217: out<=0;
   32218: out<=1;
   32219: out<=1;
   32220: out<=0;
   32221: out<=1;
   32222: out<=0;
   32223: out<=1;
   32224: out<=0;
   32225: out<=1;
   32226: out<=1;
   32227: out<=0;
   32228: out<=0;
   32229: out<=0;
   32230: out<=0;
   32231: out<=0;
   32232: out<=1;
   32233: out<=1;
   32234: out<=0;
   32235: out<=0;
   32236: out<=1;
   32237: out<=0;
   32238: out<=1;
   32239: out<=0;
   32240: out<=1;
   32241: out<=0;
   32242: out<=0;
   32243: out<=1;
   32244: out<=1;
   32245: out<=1;
   32246: out<=1;
   32247: out<=1;
   32248: out<=0;
   32249: out<=0;
   32250: out<=1;
   32251: out<=1;
   32252: out<=0;
   32253: out<=1;
   32254: out<=0;
   32255: out<=1;
   32256: out<=1;
   32257: out<=0;
   32258: out<=1;
   32259: out<=0;
   32260: out<=1;
   32261: out<=1;
   32262: out<=0;
   32263: out<=0;
   32264: out<=1;
   32265: out<=1;
   32266: out<=1;
   32267: out<=1;
   32268: out<=1;
   32269: out<=0;
   32270: out<=0;
   32271: out<=1;
   32272: out<=0;
   32273: out<=1;
   32274: out<=0;
   32275: out<=1;
   32276: out<=0;
   32277: out<=0;
   32278: out<=1;
   32279: out<=1;
   32280: out<=0;
   32281: out<=0;
   32282: out<=0;
   32283: out<=0;
   32284: out<=0;
   32285: out<=1;
   32286: out<=1;
   32287: out<=0;
   32288: out<=1;
   32289: out<=0;
   32290: out<=1;
   32291: out<=0;
   32292: out<=1;
   32293: out<=1;
   32294: out<=0;
   32295: out<=0;
   32296: out<=1;
   32297: out<=1;
   32298: out<=1;
   32299: out<=1;
   32300: out<=1;
   32301: out<=0;
   32302: out<=0;
   32303: out<=1;
   32304: out<=0;
   32305: out<=1;
   32306: out<=0;
   32307: out<=1;
   32308: out<=0;
   32309: out<=0;
   32310: out<=1;
   32311: out<=1;
   32312: out<=0;
   32313: out<=0;
   32314: out<=0;
   32315: out<=0;
   32316: out<=0;
   32317: out<=1;
   32318: out<=1;
   32319: out<=0;
   32320: out<=0;
   32321: out<=1;
   32322: out<=0;
   32323: out<=1;
   32324: out<=0;
   32325: out<=0;
   32326: out<=1;
   32327: out<=1;
   32328: out<=0;
   32329: out<=0;
   32330: out<=0;
   32331: out<=0;
   32332: out<=0;
   32333: out<=1;
   32334: out<=1;
   32335: out<=0;
   32336: out<=0;
   32337: out<=1;
   32338: out<=0;
   32339: out<=1;
   32340: out<=0;
   32341: out<=0;
   32342: out<=1;
   32343: out<=1;
   32344: out<=0;
   32345: out<=0;
   32346: out<=0;
   32347: out<=0;
   32348: out<=0;
   32349: out<=1;
   32350: out<=1;
   32351: out<=0;
   32352: out<=1;
   32353: out<=0;
   32354: out<=1;
   32355: out<=0;
   32356: out<=1;
   32357: out<=1;
   32358: out<=0;
   32359: out<=0;
   32360: out<=1;
   32361: out<=1;
   32362: out<=1;
   32363: out<=1;
   32364: out<=1;
   32365: out<=0;
   32366: out<=0;
   32367: out<=1;
   32368: out<=1;
   32369: out<=0;
   32370: out<=1;
   32371: out<=0;
   32372: out<=1;
   32373: out<=1;
   32374: out<=0;
   32375: out<=0;
   32376: out<=1;
   32377: out<=1;
   32378: out<=1;
   32379: out<=1;
   32380: out<=1;
   32381: out<=0;
   32382: out<=0;
   32383: out<=1;
   32384: out<=0;
   32385: out<=1;
   32386: out<=0;
   32387: out<=1;
   32388: out<=0;
   32389: out<=0;
   32390: out<=1;
   32391: out<=1;
   32392: out<=0;
   32393: out<=0;
   32394: out<=0;
   32395: out<=0;
   32396: out<=0;
   32397: out<=1;
   32398: out<=1;
   32399: out<=0;
   32400: out<=0;
   32401: out<=1;
   32402: out<=0;
   32403: out<=1;
   32404: out<=0;
   32405: out<=0;
   32406: out<=1;
   32407: out<=1;
   32408: out<=0;
   32409: out<=0;
   32410: out<=0;
   32411: out<=0;
   32412: out<=0;
   32413: out<=1;
   32414: out<=1;
   32415: out<=0;
   32416: out<=0;
   32417: out<=1;
   32418: out<=0;
   32419: out<=1;
   32420: out<=0;
   32421: out<=0;
   32422: out<=1;
   32423: out<=1;
   32424: out<=0;
   32425: out<=0;
   32426: out<=0;
   32427: out<=0;
   32428: out<=0;
   32429: out<=1;
   32430: out<=1;
   32431: out<=0;
   32432: out<=0;
   32433: out<=1;
   32434: out<=0;
   32435: out<=1;
   32436: out<=0;
   32437: out<=0;
   32438: out<=1;
   32439: out<=1;
   32440: out<=0;
   32441: out<=0;
   32442: out<=0;
   32443: out<=0;
   32444: out<=0;
   32445: out<=1;
   32446: out<=1;
   32447: out<=0;
   32448: out<=1;
   32449: out<=0;
   32450: out<=1;
   32451: out<=0;
   32452: out<=1;
   32453: out<=1;
   32454: out<=0;
   32455: out<=0;
   32456: out<=1;
   32457: out<=1;
   32458: out<=1;
   32459: out<=1;
   32460: out<=1;
   32461: out<=0;
   32462: out<=0;
   32463: out<=1;
   32464: out<=0;
   32465: out<=1;
   32466: out<=0;
   32467: out<=1;
   32468: out<=0;
   32469: out<=0;
   32470: out<=1;
   32471: out<=1;
   32472: out<=0;
   32473: out<=0;
   32474: out<=0;
   32475: out<=0;
   32476: out<=0;
   32477: out<=1;
   32478: out<=1;
   32479: out<=0;
   32480: out<=0;
   32481: out<=1;
   32482: out<=0;
   32483: out<=1;
   32484: out<=0;
   32485: out<=0;
   32486: out<=1;
   32487: out<=1;
   32488: out<=0;
   32489: out<=0;
   32490: out<=0;
   32491: out<=0;
   32492: out<=0;
   32493: out<=1;
   32494: out<=1;
   32495: out<=0;
   32496: out<=1;
   32497: out<=0;
   32498: out<=1;
   32499: out<=0;
   32500: out<=1;
   32501: out<=1;
   32502: out<=0;
   32503: out<=0;
   32504: out<=1;
   32505: out<=1;
   32506: out<=1;
   32507: out<=1;
   32508: out<=1;
   32509: out<=0;
   32510: out<=0;
   32511: out<=1;
   32512: out<=1;
   32513: out<=1;
   32514: out<=0;
   32515: out<=0;
   32516: out<=0;
   32517: out<=1;
   32518: out<=0;
   32519: out<=1;
   32520: out<=0;
   32521: out<=1;
   32522: out<=1;
   32523: out<=0;
   32524: out<=1;
   32525: out<=1;
   32526: out<=1;
   32527: out<=1;
   32528: out<=1;
   32529: out<=1;
   32530: out<=0;
   32531: out<=0;
   32532: out<=0;
   32533: out<=1;
   32534: out<=0;
   32535: out<=1;
   32536: out<=0;
   32537: out<=1;
   32538: out<=1;
   32539: out<=0;
   32540: out<=1;
   32541: out<=1;
   32542: out<=1;
   32543: out<=1;
   32544: out<=0;
   32545: out<=0;
   32546: out<=1;
   32547: out<=1;
   32548: out<=1;
   32549: out<=0;
   32550: out<=1;
   32551: out<=0;
   32552: out<=1;
   32553: out<=0;
   32554: out<=0;
   32555: out<=1;
   32556: out<=0;
   32557: out<=0;
   32558: out<=0;
   32559: out<=0;
   32560: out<=0;
   32561: out<=0;
   32562: out<=1;
   32563: out<=1;
   32564: out<=1;
   32565: out<=0;
   32566: out<=1;
   32567: out<=0;
   32568: out<=1;
   32569: out<=0;
   32570: out<=0;
   32571: out<=1;
   32572: out<=0;
   32573: out<=0;
   32574: out<=0;
   32575: out<=0;
   32576: out<=0;
   32577: out<=0;
   32578: out<=1;
   32579: out<=1;
   32580: out<=1;
   32581: out<=0;
   32582: out<=1;
   32583: out<=0;
   32584: out<=1;
   32585: out<=0;
   32586: out<=0;
   32587: out<=1;
   32588: out<=0;
   32589: out<=0;
   32590: out<=0;
   32591: out<=0;
   32592: out<=1;
   32593: out<=1;
   32594: out<=0;
   32595: out<=0;
   32596: out<=0;
   32597: out<=1;
   32598: out<=0;
   32599: out<=1;
   32600: out<=0;
   32601: out<=1;
   32602: out<=1;
   32603: out<=0;
   32604: out<=1;
   32605: out<=1;
   32606: out<=1;
   32607: out<=1;
   32608: out<=0;
   32609: out<=0;
   32610: out<=1;
   32611: out<=1;
   32612: out<=1;
   32613: out<=0;
   32614: out<=1;
   32615: out<=0;
   32616: out<=1;
   32617: out<=0;
   32618: out<=0;
   32619: out<=1;
   32620: out<=0;
   32621: out<=0;
   32622: out<=0;
   32623: out<=0;
   32624: out<=1;
   32625: out<=1;
   32626: out<=0;
   32627: out<=0;
   32628: out<=0;
   32629: out<=1;
   32630: out<=0;
   32631: out<=1;
   32632: out<=0;
   32633: out<=1;
   32634: out<=1;
   32635: out<=0;
   32636: out<=1;
   32637: out<=1;
   32638: out<=1;
   32639: out<=1;
   32640: out<=0;
   32641: out<=0;
   32642: out<=1;
   32643: out<=1;
   32644: out<=1;
   32645: out<=0;
   32646: out<=1;
   32647: out<=0;
   32648: out<=1;
   32649: out<=0;
   32650: out<=0;
   32651: out<=1;
   32652: out<=0;
   32653: out<=0;
   32654: out<=0;
   32655: out<=0;
   32656: out<=1;
   32657: out<=1;
   32658: out<=0;
   32659: out<=0;
   32660: out<=0;
   32661: out<=1;
   32662: out<=0;
   32663: out<=1;
   32664: out<=0;
   32665: out<=1;
   32666: out<=1;
   32667: out<=0;
   32668: out<=1;
   32669: out<=1;
   32670: out<=1;
   32671: out<=1;
   32672: out<=1;
   32673: out<=1;
   32674: out<=0;
   32675: out<=0;
   32676: out<=0;
   32677: out<=1;
   32678: out<=0;
   32679: out<=1;
   32680: out<=0;
   32681: out<=1;
   32682: out<=1;
   32683: out<=0;
   32684: out<=1;
   32685: out<=1;
   32686: out<=1;
   32687: out<=1;
   32688: out<=0;
   32689: out<=0;
   32690: out<=1;
   32691: out<=1;
   32692: out<=1;
   32693: out<=0;
   32694: out<=1;
   32695: out<=0;
   32696: out<=1;
   32697: out<=0;
   32698: out<=0;
   32699: out<=1;
   32700: out<=0;
   32701: out<=0;
   32702: out<=0;
   32703: out<=0;
   32704: out<=1;
   32705: out<=1;
   32706: out<=0;
   32707: out<=0;
   32708: out<=0;
   32709: out<=1;
   32710: out<=0;
   32711: out<=1;
   32712: out<=0;
   32713: out<=1;
   32714: out<=1;
   32715: out<=0;
   32716: out<=1;
   32717: out<=1;
   32718: out<=1;
   32719: out<=1;
   32720: out<=1;
   32721: out<=1;
   32722: out<=0;
   32723: out<=0;
   32724: out<=0;
   32725: out<=1;
   32726: out<=0;
   32727: out<=1;
   32728: out<=0;
   32729: out<=1;
   32730: out<=1;
   32731: out<=0;
   32732: out<=1;
   32733: out<=1;
   32734: out<=1;
   32735: out<=1;
   32736: out<=1;
   32737: out<=1;
   32738: out<=0;
   32739: out<=0;
   32740: out<=0;
   32741: out<=1;
   32742: out<=0;
   32743: out<=1;
   32744: out<=0;
   32745: out<=1;
   32746: out<=1;
   32747: out<=0;
   32748: out<=1;
   32749: out<=1;
   32750: out<=1;
   32751: out<=1;
   32752: out<=1;
   32753: out<=1;
   32754: out<=0;
   32755: out<=0;
   32756: out<=0;
   32757: out<=1;
   32758: out<=0;
   32759: out<=1;
   32760: out<=0;
   32761: out<=1;
   32762: out<=1;
   32763: out<=0;
   32764: out<=1;
   32765: out<=1;
   32766: out<=1;
   32767: out<=1;
   32768: out<=0;
   32769: out<=0;
   32770: out<=0;
   32771: out<=0;
   32772: out<=1;
   32773: out<=0;
   32774: out<=0;
   32775: out<=1;
   32776: out<=0;
   32777: out<=1;
   32778: out<=0;
   32779: out<=1;
   32780: out<=1;
   32781: out<=1;
   32782: out<=0;
   32783: out<=0;
   32784: out<=0;
   32785: out<=0;
   32786: out<=0;
   32787: out<=0;
   32788: out<=1;
   32789: out<=0;
   32790: out<=0;
   32791: out<=1;
   32792: out<=0;
   32793: out<=1;
   32794: out<=0;
   32795: out<=1;
   32796: out<=1;
   32797: out<=1;
   32798: out<=0;
   32799: out<=0;
   32800: out<=0;
   32801: out<=0;
   32802: out<=0;
   32803: out<=0;
   32804: out<=1;
   32805: out<=0;
   32806: out<=0;
   32807: out<=1;
   32808: out<=0;
   32809: out<=1;
   32810: out<=0;
   32811: out<=1;
   32812: out<=1;
   32813: out<=1;
   32814: out<=0;
   32815: out<=0;
   32816: out<=0;
   32817: out<=0;
   32818: out<=0;
   32819: out<=0;
   32820: out<=1;
   32821: out<=0;
   32822: out<=0;
   32823: out<=1;
   32824: out<=0;
   32825: out<=1;
   32826: out<=0;
   32827: out<=1;
   32828: out<=1;
   32829: out<=1;
   32830: out<=0;
   32831: out<=0;
   32832: out<=1;
   32833: out<=1;
   32834: out<=1;
   32835: out<=1;
   32836: out<=0;
   32837: out<=1;
   32838: out<=1;
   32839: out<=0;
   32840: out<=1;
   32841: out<=0;
   32842: out<=1;
   32843: out<=0;
   32844: out<=0;
   32845: out<=0;
   32846: out<=1;
   32847: out<=1;
   32848: out<=0;
   32849: out<=0;
   32850: out<=0;
   32851: out<=0;
   32852: out<=1;
   32853: out<=0;
   32854: out<=0;
   32855: out<=1;
   32856: out<=0;
   32857: out<=1;
   32858: out<=0;
   32859: out<=1;
   32860: out<=1;
   32861: out<=1;
   32862: out<=0;
   32863: out<=0;
   32864: out<=0;
   32865: out<=0;
   32866: out<=0;
   32867: out<=0;
   32868: out<=1;
   32869: out<=0;
   32870: out<=0;
   32871: out<=1;
   32872: out<=0;
   32873: out<=1;
   32874: out<=0;
   32875: out<=1;
   32876: out<=1;
   32877: out<=1;
   32878: out<=0;
   32879: out<=0;
   32880: out<=1;
   32881: out<=1;
   32882: out<=1;
   32883: out<=1;
   32884: out<=0;
   32885: out<=1;
   32886: out<=1;
   32887: out<=0;
   32888: out<=1;
   32889: out<=0;
   32890: out<=1;
   32891: out<=0;
   32892: out<=0;
   32893: out<=0;
   32894: out<=1;
   32895: out<=1;
   32896: out<=0;
   32897: out<=0;
   32898: out<=0;
   32899: out<=0;
   32900: out<=1;
   32901: out<=0;
   32902: out<=0;
   32903: out<=1;
   32904: out<=0;
   32905: out<=1;
   32906: out<=0;
   32907: out<=1;
   32908: out<=1;
   32909: out<=1;
   32910: out<=0;
   32911: out<=0;
   32912: out<=1;
   32913: out<=1;
   32914: out<=1;
   32915: out<=1;
   32916: out<=0;
   32917: out<=1;
   32918: out<=1;
   32919: out<=0;
   32920: out<=1;
   32921: out<=0;
   32922: out<=1;
   32923: out<=0;
   32924: out<=0;
   32925: out<=0;
   32926: out<=1;
   32927: out<=1;
   32928: out<=0;
   32929: out<=0;
   32930: out<=0;
   32931: out<=0;
   32932: out<=1;
   32933: out<=0;
   32934: out<=0;
   32935: out<=1;
   32936: out<=0;
   32937: out<=1;
   32938: out<=0;
   32939: out<=1;
   32940: out<=1;
   32941: out<=1;
   32942: out<=0;
   32943: out<=0;
   32944: out<=1;
   32945: out<=1;
   32946: out<=1;
   32947: out<=1;
   32948: out<=0;
   32949: out<=1;
   32950: out<=1;
   32951: out<=0;
   32952: out<=1;
   32953: out<=0;
   32954: out<=1;
   32955: out<=0;
   32956: out<=0;
   32957: out<=0;
   32958: out<=1;
   32959: out<=1;
   32960: out<=1;
   32961: out<=1;
   32962: out<=1;
   32963: out<=1;
   32964: out<=0;
   32965: out<=1;
   32966: out<=1;
   32967: out<=0;
   32968: out<=1;
   32969: out<=0;
   32970: out<=1;
   32971: out<=0;
   32972: out<=0;
   32973: out<=0;
   32974: out<=1;
   32975: out<=1;
   32976: out<=1;
   32977: out<=1;
   32978: out<=1;
   32979: out<=1;
   32980: out<=0;
   32981: out<=1;
   32982: out<=1;
   32983: out<=0;
   32984: out<=1;
   32985: out<=0;
   32986: out<=1;
   32987: out<=0;
   32988: out<=0;
   32989: out<=0;
   32990: out<=1;
   32991: out<=1;
   32992: out<=0;
   32993: out<=0;
   32994: out<=0;
   32995: out<=0;
   32996: out<=1;
   32997: out<=0;
   32998: out<=0;
   32999: out<=1;
   33000: out<=0;
   33001: out<=1;
   33002: out<=0;
   33003: out<=1;
   33004: out<=1;
   33005: out<=1;
   33006: out<=0;
   33007: out<=0;
   33008: out<=0;
   33009: out<=0;
   33010: out<=0;
   33011: out<=0;
   33012: out<=1;
   33013: out<=0;
   33014: out<=0;
   33015: out<=1;
   33016: out<=0;
   33017: out<=1;
   33018: out<=0;
   33019: out<=1;
   33020: out<=1;
   33021: out<=1;
   33022: out<=0;
   33023: out<=0;
   33024: out<=0;
   33025: out<=1;
   33026: out<=1;
   33027: out<=0;
   33028: out<=0;
   33029: out<=0;
   33030: out<=0;
   33031: out<=0;
   33032: out<=1;
   33033: out<=1;
   33034: out<=0;
   33035: out<=0;
   33036: out<=1;
   33037: out<=0;
   33038: out<=1;
   33039: out<=0;
   33040: out<=1;
   33041: out<=0;
   33042: out<=0;
   33043: out<=1;
   33044: out<=1;
   33045: out<=1;
   33046: out<=1;
   33047: out<=1;
   33048: out<=0;
   33049: out<=0;
   33050: out<=1;
   33051: out<=1;
   33052: out<=0;
   33053: out<=1;
   33054: out<=0;
   33055: out<=1;
   33056: out<=1;
   33057: out<=0;
   33058: out<=0;
   33059: out<=1;
   33060: out<=1;
   33061: out<=1;
   33062: out<=1;
   33063: out<=1;
   33064: out<=0;
   33065: out<=0;
   33066: out<=1;
   33067: out<=1;
   33068: out<=0;
   33069: out<=1;
   33070: out<=0;
   33071: out<=1;
   33072: out<=0;
   33073: out<=1;
   33074: out<=1;
   33075: out<=0;
   33076: out<=0;
   33077: out<=0;
   33078: out<=0;
   33079: out<=0;
   33080: out<=1;
   33081: out<=1;
   33082: out<=0;
   33083: out<=0;
   33084: out<=1;
   33085: out<=0;
   33086: out<=1;
   33087: out<=0;
   33088: out<=1;
   33089: out<=0;
   33090: out<=0;
   33091: out<=1;
   33092: out<=1;
   33093: out<=1;
   33094: out<=1;
   33095: out<=1;
   33096: out<=0;
   33097: out<=0;
   33098: out<=1;
   33099: out<=1;
   33100: out<=0;
   33101: out<=1;
   33102: out<=0;
   33103: out<=1;
   33104: out<=1;
   33105: out<=0;
   33106: out<=0;
   33107: out<=1;
   33108: out<=1;
   33109: out<=1;
   33110: out<=1;
   33111: out<=1;
   33112: out<=0;
   33113: out<=0;
   33114: out<=1;
   33115: out<=1;
   33116: out<=0;
   33117: out<=1;
   33118: out<=0;
   33119: out<=1;
   33120: out<=1;
   33121: out<=0;
   33122: out<=0;
   33123: out<=1;
   33124: out<=1;
   33125: out<=1;
   33126: out<=1;
   33127: out<=1;
   33128: out<=0;
   33129: out<=0;
   33130: out<=1;
   33131: out<=1;
   33132: out<=0;
   33133: out<=1;
   33134: out<=0;
   33135: out<=1;
   33136: out<=1;
   33137: out<=0;
   33138: out<=0;
   33139: out<=1;
   33140: out<=1;
   33141: out<=1;
   33142: out<=1;
   33143: out<=1;
   33144: out<=0;
   33145: out<=0;
   33146: out<=1;
   33147: out<=1;
   33148: out<=0;
   33149: out<=1;
   33150: out<=0;
   33151: out<=1;
   33152: out<=0;
   33153: out<=1;
   33154: out<=1;
   33155: out<=0;
   33156: out<=0;
   33157: out<=0;
   33158: out<=0;
   33159: out<=0;
   33160: out<=1;
   33161: out<=1;
   33162: out<=0;
   33163: out<=0;
   33164: out<=1;
   33165: out<=0;
   33166: out<=1;
   33167: out<=0;
   33168: out<=0;
   33169: out<=1;
   33170: out<=1;
   33171: out<=0;
   33172: out<=0;
   33173: out<=0;
   33174: out<=0;
   33175: out<=0;
   33176: out<=1;
   33177: out<=1;
   33178: out<=0;
   33179: out<=0;
   33180: out<=1;
   33181: out<=0;
   33182: out<=1;
   33183: out<=0;
   33184: out<=1;
   33185: out<=0;
   33186: out<=0;
   33187: out<=1;
   33188: out<=1;
   33189: out<=1;
   33190: out<=1;
   33191: out<=1;
   33192: out<=0;
   33193: out<=0;
   33194: out<=1;
   33195: out<=1;
   33196: out<=0;
   33197: out<=1;
   33198: out<=0;
   33199: out<=1;
   33200: out<=1;
   33201: out<=0;
   33202: out<=0;
   33203: out<=1;
   33204: out<=1;
   33205: out<=1;
   33206: out<=1;
   33207: out<=1;
   33208: out<=0;
   33209: out<=0;
   33210: out<=1;
   33211: out<=1;
   33212: out<=0;
   33213: out<=1;
   33214: out<=0;
   33215: out<=1;
   33216: out<=1;
   33217: out<=0;
   33218: out<=0;
   33219: out<=1;
   33220: out<=1;
   33221: out<=1;
   33222: out<=1;
   33223: out<=1;
   33224: out<=0;
   33225: out<=0;
   33226: out<=1;
   33227: out<=1;
   33228: out<=0;
   33229: out<=1;
   33230: out<=0;
   33231: out<=1;
   33232: out<=0;
   33233: out<=1;
   33234: out<=1;
   33235: out<=0;
   33236: out<=0;
   33237: out<=0;
   33238: out<=0;
   33239: out<=0;
   33240: out<=1;
   33241: out<=1;
   33242: out<=0;
   33243: out<=0;
   33244: out<=1;
   33245: out<=0;
   33246: out<=1;
   33247: out<=0;
   33248: out<=1;
   33249: out<=0;
   33250: out<=0;
   33251: out<=1;
   33252: out<=1;
   33253: out<=1;
   33254: out<=1;
   33255: out<=1;
   33256: out<=0;
   33257: out<=0;
   33258: out<=1;
   33259: out<=1;
   33260: out<=0;
   33261: out<=1;
   33262: out<=0;
   33263: out<=1;
   33264: out<=0;
   33265: out<=1;
   33266: out<=1;
   33267: out<=0;
   33268: out<=0;
   33269: out<=0;
   33270: out<=0;
   33271: out<=0;
   33272: out<=1;
   33273: out<=1;
   33274: out<=0;
   33275: out<=0;
   33276: out<=1;
   33277: out<=0;
   33278: out<=1;
   33279: out<=0;
   33280: out<=0;
   33281: out<=1;
   33282: out<=0;
   33283: out<=1;
   33284: out<=0;
   33285: out<=0;
   33286: out<=1;
   33287: out<=1;
   33288: out<=0;
   33289: out<=0;
   33290: out<=0;
   33291: out<=0;
   33292: out<=0;
   33293: out<=1;
   33294: out<=1;
   33295: out<=0;
   33296: out<=1;
   33297: out<=0;
   33298: out<=1;
   33299: out<=0;
   33300: out<=1;
   33301: out<=1;
   33302: out<=0;
   33303: out<=0;
   33304: out<=1;
   33305: out<=1;
   33306: out<=1;
   33307: out<=1;
   33308: out<=1;
   33309: out<=0;
   33310: out<=0;
   33311: out<=1;
   33312: out<=0;
   33313: out<=1;
   33314: out<=0;
   33315: out<=1;
   33316: out<=0;
   33317: out<=0;
   33318: out<=1;
   33319: out<=1;
   33320: out<=0;
   33321: out<=0;
   33322: out<=0;
   33323: out<=0;
   33324: out<=0;
   33325: out<=1;
   33326: out<=1;
   33327: out<=0;
   33328: out<=1;
   33329: out<=0;
   33330: out<=1;
   33331: out<=0;
   33332: out<=1;
   33333: out<=1;
   33334: out<=0;
   33335: out<=0;
   33336: out<=1;
   33337: out<=1;
   33338: out<=1;
   33339: out<=1;
   33340: out<=1;
   33341: out<=0;
   33342: out<=0;
   33343: out<=1;
   33344: out<=1;
   33345: out<=0;
   33346: out<=1;
   33347: out<=0;
   33348: out<=1;
   33349: out<=1;
   33350: out<=0;
   33351: out<=0;
   33352: out<=1;
   33353: out<=1;
   33354: out<=1;
   33355: out<=1;
   33356: out<=1;
   33357: out<=0;
   33358: out<=0;
   33359: out<=1;
   33360: out<=1;
   33361: out<=0;
   33362: out<=1;
   33363: out<=0;
   33364: out<=1;
   33365: out<=1;
   33366: out<=0;
   33367: out<=0;
   33368: out<=1;
   33369: out<=1;
   33370: out<=1;
   33371: out<=1;
   33372: out<=1;
   33373: out<=0;
   33374: out<=0;
   33375: out<=1;
   33376: out<=0;
   33377: out<=1;
   33378: out<=0;
   33379: out<=1;
   33380: out<=0;
   33381: out<=0;
   33382: out<=1;
   33383: out<=1;
   33384: out<=0;
   33385: out<=0;
   33386: out<=0;
   33387: out<=0;
   33388: out<=0;
   33389: out<=1;
   33390: out<=1;
   33391: out<=0;
   33392: out<=0;
   33393: out<=1;
   33394: out<=0;
   33395: out<=1;
   33396: out<=0;
   33397: out<=0;
   33398: out<=1;
   33399: out<=1;
   33400: out<=0;
   33401: out<=0;
   33402: out<=0;
   33403: out<=0;
   33404: out<=0;
   33405: out<=1;
   33406: out<=1;
   33407: out<=0;
   33408: out<=0;
   33409: out<=1;
   33410: out<=0;
   33411: out<=1;
   33412: out<=0;
   33413: out<=0;
   33414: out<=1;
   33415: out<=1;
   33416: out<=0;
   33417: out<=0;
   33418: out<=0;
   33419: out<=0;
   33420: out<=0;
   33421: out<=1;
   33422: out<=1;
   33423: out<=0;
   33424: out<=0;
   33425: out<=1;
   33426: out<=0;
   33427: out<=1;
   33428: out<=0;
   33429: out<=0;
   33430: out<=1;
   33431: out<=1;
   33432: out<=0;
   33433: out<=0;
   33434: out<=0;
   33435: out<=0;
   33436: out<=0;
   33437: out<=1;
   33438: out<=1;
   33439: out<=0;
   33440: out<=0;
   33441: out<=1;
   33442: out<=0;
   33443: out<=1;
   33444: out<=0;
   33445: out<=0;
   33446: out<=1;
   33447: out<=1;
   33448: out<=0;
   33449: out<=0;
   33450: out<=0;
   33451: out<=0;
   33452: out<=0;
   33453: out<=1;
   33454: out<=1;
   33455: out<=0;
   33456: out<=0;
   33457: out<=1;
   33458: out<=0;
   33459: out<=1;
   33460: out<=0;
   33461: out<=0;
   33462: out<=1;
   33463: out<=1;
   33464: out<=0;
   33465: out<=0;
   33466: out<=0;
   33467: out<=0;
   33468: out<=0;
   33469: out<=1;
   33470: out<=1;
   33471: out<=0;
   33472: out<=1;
   33473: out<=0;
   33474: out<=1;
   33475: out<=0;
   33476: out<=1;
   33477: out<=1;
   33478: out<=0;
   33479: out<=0;
   33480: out<=1;
   33481: out<=1;
   33482: out<=1;
   33483: out<=1;
   33484: out<=1;
   33485: out<=0;
   33486: out<=0;
   33487: out<=1;
   33488: out<=0;
   33489: out<=1;
   33490: out<=0;
   33491: out<=1;
   33492: out<=0;
   33493: out<=0;
   33494: out<=1;
   33495: out<=1;
   33496: out<=0;
   33497: out<=0;
   33498: out<=0;
   33499: out<=0;
   33500: out<=0;
   33501: out<=1;
   33502: out<=1;
   33503: out<=0;
   33504: out<=0;
   33505: out<=1;
   33506: out<=0;
   33507: out<=1;
   33508: out<=0;
   33509: out<=0;
   33510: out<=1;
   33511: out<=1;
   33512: out<=0;
   33513: out<=0;
   33514: out<=0;
   33515: out<=0;
   33516: out<=0;
   33517: out<=1;
   33518: out<=1;
   33519: out<=0;
   33520: out<=1;
   33521: out<=0;
   33522: out<=1;
   33523: out<=0;
   33524: out<=1;
   33525: out<=1;
   33526: out<=0;
   33527: out<=0;
   33528: out<=1;
   33529: out<=1;
   33530: out<=1;
   33531: out<=1;
   33532: out<=1;
   33533: out<=0;
   33534: out<=0;
   33535: out<=1;
   33536: out<=0;
   33537: out<=0;
   33538: out<=1;
   33539: out<=1;
   33540: out<=1;
   33541: out<=0;
   33542: out<=1;
   33543: out<=0;
   33544: out<=1;
   33545: out<=0;
   33546: out<=0;
   33547: out<=1;
   33548: out<=0;
   33549: out<=0;
   33550: out<=0;
   33551: out<=0;
   33552: out<=0;
   33553: out<=0;
   33554: out<=1;
   33555: out<=1;
   33556: out<=1;
   33557: out<=0;
   33558: out<=1;
   33559: out<=0;
   33560: out<=1;
   33561: out<=0;
   33562: out<=0;
   33563: out<=1;
   33564: out<=0;
   33565: out<=0;
   33566: out<=0;
   33567: out<=0;
   33568: out<=1;
   33569: out<=1;
   33570: out<=0;
   33571: out<=0;
   33572: out<=0;
   33573: out<=1;
   33574: out<=0;
   33575: out<=1;
   33576: out<=0;
   33577: out<=1;
   33578: out<=1;
   33579: out<=0;
   33580: out<=1;
   33581: out<=1;
   33582: out<=1;
   33583: out<=1;
   33584: out<=1;
   33585: out<=1;
   33586: out<=0;
   33587: out<=0;
   33588: out<=0;
   33589: out<=1;
   33590: out<=0;
   33591: out<=1;
   33592: out<=0;
   33593: out<=1;
   33594: out<=1;
   33595: out<=0;
   33596: out<=1;
   33597: out<=1;
   33598: out<=1;
   33599: out<=1;
   33600: out<=1;
   33601: out<=1;
   33602: out<=0;
   33603: out<=0;
   33604: out<=0;
   33605: out<=1;
   33606: out<=0;
   33607: out<=1;
   33608: out<=0;
   33609: out<=1;
   33610: out<=1;
   33611: out<=0;
   33612: out<=1;
   33613: out<=1;
   33614: out<=1;
   33615: out<=1;
   33616: out<=0;
   33617: out<=0;
   33618: out<=1;
   33619: out<=1;
   33620: out<=1;
   33621: out<=0;
   33622: out<=1;
   33623: out<=0;
   33624: out<=1;
   33625: out<=0;
   33626: out<=0;
   33627: out<=1;
   33628: out<=0;
   33629: out<=0;
   33630: out<=0;
   33631: out<=0;
   33632: out<=1;
   33633: out<=1;
   33634: out<=0;
   33635: out<=0;
   33636: out<=0;
   33637: out<=1;
   33638: out<=0;
   33639: out<=1;
   33640: out<=0;
   33641: out<=1;
   33642: out<=1;
   33643: out<=0;
   33644: out<=1;
   33645: out<=1;
   33646: out<=1;
   33647: out<=1;
   33648: out<=0;
   33649: out<=0;
   33650: out<=1;
   33651: out<=1;
   33652: out<=1;
   33653: out<=0;
   33654: out<=1;
   33655: out<=0;
   33656: out<=1;
   33657: out<=0;
   33658: out<=0;
   33659: out<=1;
   33660: out<=0;
   33661: out<=0;
   33662: out<=0;
   33663: out<=0;
   33664: out<=0;
   33665: out<=0;
   33666: out<=1;
   33667: out<=1;
   33668: out<=1;
   33669: out<=0;
   33670: out<=1;
   33671: out<=0;
   33672: out<=1;
   33673: out<=0;
   33674: out<=0;
   33675: out<=1;
   33676: out<=0;
   33677: out<=0;
   33678: out<=0;
   33679: out<=0;
   33680: out<=1;
   33681: out<=1;
   33682: out<=0;
   33683: out<=0;
   33684: out<=0;
   33685: out<=1;
   33686: out<=0;
   33687: out<=1;
   33688: out<=0;
   33689: out<=1;
   33690: out<=1;
   33691: out<=0;
   33692: out<=1;
   33693: out<=1;
   33694: out<=1;
   33695: out<=1;
   33696: out<=1;
   33697: out<=1;
   33698: out<=0;
   33699: out<=0;
   33700: out<=0;
   33701: out<=1;
   33702: out<=0;
   33703: out<=1;
   33704: out<=0;
   33705: out<=1;
   33706: out<=1;
   33707: out<=0;
   33708: out<=1;
   33709: out<=1;
   33710: out<=1;
   33711: out<=1;
   33712: out<=0;
   33713: out<=0;
   33714: out<=1;
   33715: out<=1;
   33716: out<=1;
   33717: out<=0;
   33718: out<=1;
   33719: out<=0;
   33720: out<=1;
   33721: out<=0;
   33722: out<=0;
   33723: out<=1;
   33724: out<=0;
   33725: out<=0;
   33726: out<=0;
   33727: out<=0;
   33728: out<=1;
   33729: out<=1;
   33730: out<=0;
   33731: out<=0;
   33732: out<=0;
   33733: out<=1;
   33734: out<=0;
   33735: out<=1;
   33736: out<=0;
   33737: out<=1;
   33738: out<=1;
   33739: out<=0;
   33740: out<=1;
   33741: out<=1;
   33742: out<=1;
   33743: out<=1;
   33744: out<=1;
   33745: out<=1;
   33746: out<=0;
   33747: out<=0;
   33748: out<=0;
   33749: out<=1;
   33750: out<=0;
   33751: out<=1;
   33752: out<=0;
   33753: out<=1;
   33754: out<=1;
   33755: out<=0;
   33756: out<=1;
   33757: out<=1;
   33758: out<=1;
   33759: out<=1;
   33760: out<=1;
   33761: out<=1;
   33762: out<=0;
   33763: out<=0;
   33764: out<=0;
   33765: out<=1;
   33766: out<=0;
   33767: out<=1;
   33768: out<=0;
   33769: out<=1;
   33770: out<=1;
   33771: out<=0;
   33772: out<=1;
   33773: out<=1;
   33774: out<=1;
   33775: out<=1;
   33776: out<=1;
   33777: out<=1;
   33778: out<=0;
   33779: out<=0;
   33780: out<=0;
   33781: out<=1;
   33782: out<=0;
   33783: out<=1;
   33784: out<=0;
   33785: out<=1;
   33786: out<=1;
   33787: out<=0;
   33788: out<=1;
   33789: out<=1;
   33790: out<=1;
   33791: out<=1;
   33792: out<=0;
   33793: out<=1;
   33794: out<=1;
   33795: out<=0;
   33796: out<=1;
   33797: out<=1;
   33798: out<=1;
   33799: out<=1;
   33800: out<=0;
   33801: out<=0;
   33802: out<=1;
   33803: out<=1;
   33804: out<=1;
   33805: out<=0;
   33806: out<=1;
   33807: out<=0;
   33808: out<=0;
   33809: out<=1;
   33810: out<=1;
   33811: out<=0;
   33812: out<=1;
   33813: out<=1;
   33814: out<=1;
   33815: out<=1;
   33816: out<=0;
   33817: out<=0;
   33818: out<=1;
   33819: out<=1;
   33820: out<=1;
   33821: out<=0;
   33822: out<=1;
   33823: out<=0;
   33824: out<=0;
   33825: out<=1;
   33826: out<=1;
   33827: out<=0;
   33828: out<=1;
   33829: out<=1;
   33830: out<=1;
   33831: out<=1;
   33832: out<=0;
   33833: out<=0;
   33834: out<=1;
   33835: out<=1;
   33836: out<=1;
   33837: out<=0;
   33838: out<=1;
   33839: out<=0;
   33840: out<=0;
   33841: out<=1;
   33842: out<=1;
   33843: out<=0;
   33844: out<=1;
   33845: out<=1;
   33846: out<=1;
   33847: out<=1;
   33848: out<=0;
   33849: out<=0;
   33850: out<=1;
   33851: out<=1;
   33852: out<=1;
   33853: out<=0;
   33854: out<=1;
   33855: out<=0;
   33856: out<=1;
   33857: out<=0;
   33858: out<=0;
   33859: out<=1;
   33860: out<=0;
   33861: out<=0;
   33862: out<=0;
   33863: out<=0;
   33864: out<=1;
   33865: out<=1;
   33866: out<=0;
   33867: out<=0;
   33868: out<=0;
   33869: out<=1;
   33870: out<=0;
   33871: out<=1;
   33872: out<=0;
   33873: out<=1;
   33874: out<=1;
   33875: out<=0;
   33876: out<=1;
   33877: out<=1;
   33878: out<=1;
   33879: out<=1;
   33880: out<=0;
   33881: out<=0;
   33882: out<=1;
   33883: out<=1;
   33884: out<=1;
   33885: out<=0;
   33886: out<=1;
   33887: out<=0;
   33888: out<=0;
   33889: out<=1;
   33890: out<=1;
   33891: out<=0;
   33892: out<=1;
   33893: out<=1;
   33894: out<=1;
   33895: out<=1;
   33896: out<=0;
   33897: out<=0;
   33898: out<=1;
   33899: out<=1;
   33900: out<=1;
   33901: out<=0;
   33902: out<=1;
   33903: out<=0;
   33904: out<=1;
   33905: out<=0;
   33906: out<=0;
   33907: out<=1;
   33908: out<=0;
   33909: out<=0;
   33910: out<=0;
   33911: out<=0;
   33912: out<=1;
   33913: out<=1;
   33914: out<=0;
   33915: out<=0;
   33916: out<=0;
   33917: out<=1;
   33918: out<=0;
   33919: out<=1;
   33920: out<=0;
   33921: out<=1;
   33922: out<=1;
   33923: out<=0;
   33924: out<=1;
   33925: out<=1;
   33926: out<=1;
   33927: out<=1;
   33928: out<=0;
   33929: out<=0;
   33930: out<=1;
   33931: out<=1;
   33932: out<=1;
   33933: out<=0;
   33934: out<=1;
   33935: out<=0;
   33936: out<=1;
   33937: out<=0;
   33938: out<=0;
   33939: out<=1;
   33940: out<=0;
   33941: out<=0;
   33942: out<=0;
   33943: out<=0;
   33944: out<=1;
   33945: out<=1;
   33946: out<=0;
   33947: out<=0;
   33948: out<=0;
   33949: out<=1;
   33950: out<=0;
   33951: out<=1;
   33952: out<=0;
   33953: out<=1;
   33954: out<=1;
   33955: out<=0;
   33956: out<=1;
   33957: out<=1;
   33958: out<=1;
   33959: out<=1;
   33960: out<=0;
   33961: out<=0;
   33962: out<=1;
   33963: out<=1;
   33964: out<=1;
   33965: out<=0;
   33966: out<=1;
   33967: out<=0;
   33968: out<=1;
   33969: out<=0;
   33970: out<=0;
   33971: out<=1;
   33972: out<=0;
   33973: out<=0;
   33974: out<=0;
   33975: out<=0;
   33976: out<=1;
   33977: out<=1;
   33978: out<=0;
   33979: out<=0;
   33980: out<=0;
   33981: out<=1;
   33982: out<=0;
   33983: out<=1;
   33984: out<=1;
   33985: out<=0;
   33986: out<=0;
   33987: out<=1;
   33988: out<=0;
   33989: out<=0;
   33990: out<=0;
   33991: out<=0;
   33992: out<=1;
   33993: out<=1;
   33994: out<=0;
   33995: out<=0;
   33996: out<=0;
   33997: out<=1;
   33998: out<=0;
   33999: out<=1;
   34000: out<=1;
   34001: out<=0;
   34002: out<=0;
   34003: out<=1;
   34004: out<=0;
   34005: out<=0;
   34006: out<=0;
   34007: out<=0;
   34008: out<=1;
   34009: out<=1;
   34010: out<=0;
   34011: out<=0;
   34012: out<=0;
   34013: out<=1;
   34014: out<=0;
   34015: out<=1;
   34016: out<=0;
   34017: out<=1;
   34018: out<=1;
   34019: out<=0;
   34020: out<=1;
   34021: out<=1;
   34022: out<=1;
   34023: out<=1;
   34024: out<=0;
   34025: out<=0;
   34026: out<=1;
   34027: out<=1;
   34028: out<=1;
   34029: out<=0;
   34030: out<=1;
   34031: out<=0;
   34032: out<=0;
   34033: out<=1;
   34034: out<=1;
   34035: out<=0;
   34036: out<=1;
   34037: out<=1;
   34038: out<=1;
   34039: out<=1;
   34040: out<=0;
   34041: out<=0;
   34042: out<=1;
   34043: out<=1;
   34044: out<=1;
   34045: out<=0;
   34046: out<=1;
   34047: out<=0;
   34048: out<=1;
   34049: out<=1;
   34050: out<=1;
   34051: out<=1;
   34052: out<=1;
   34053: out<=0;
   34054: out<=0;
   34055: out<=1;
   34056: out<=0;
   34057: out<=1;
   34058: out<=0;
   34059: out<=1;
   34060: out<=0;
   34061: out<=0;
   34062: out<=1;
   34063: out<=1;
   34064: out<=0;
   34065: out<=0;
   34066: out<=0;
   34067: out<=0;
   34068: out<=0;
   34069: out<=1;
   34070: out<=1;
   34071: out<=0;
   34072: out<=1;
   34073: out<=0;
   34074: out<=1;
   34075: out<=0;
   34076: out<=1;
   34077: out<=1;
   34078: out<=0;
   34079: out<=0;
   34080: out<=0;
   34081: out<=0;
   34082: out<=0;
   34083: out<=0;
   34084: out<=0;
   34085: out<=1;
   34086: out<=1;
   34087: out<=0;
   34088: out<=1;
   34089: out<=0;
   34090: out<=1;
   34091: out<=0;
   34092: out<=1;
   34093: out<=1;
   34094: out<=0;
   34095: out<=0;
   34096: out<=1;
   34097: out<=1;
   34098: out<=1;
   34099: out<=1;
   34100: out<=1;
   34101: out<=0;
   34102: out<=0;
   34103: out<=1;
   34104: out<=0;
   34105: out<=1;
   34106: out<=0;
   34107: out<=1;
   34108: out<=0;
   34109: out<=0;
   34110: out<=1;
   34111: out<=1;
   34112: out<=0;
   34113: out<=0;
   34114: out<=0;
   34115: out<=0;
   34116: out<=0;
   34117: out<=1;
   34118: out<=1;
   34119: out<=0;
   34120: out<=1;
   34121: out<=0;
   34122: out<=1;
   34123: out<=0;
   34124: out<=1;
   34125: out<=1;
   34126: out<=0;
   34127: out<=0;
   34128: out<=0;
   34129: out<=0;
   34130: out<=0;
   34131: out<=0;
   34132: out<=0;
   34133: out<=1;
   34134: out<=1;
   34135: out<=0;
   34136: out<=1;
   34137: out<=0;
   34138: out<=1;
   34139: out<=0;
   34140: out<=1;
   34141: out<=1;
   34142: out<=0;
   34143: out<=0;
   34144: out<=0;
   34145: out<=0;
   34146: out<=0;
   34147: out<=0;
   34148: out<=0;
   34149: out<=1;
   34150: out<=1;
   34151: out<=0;
   34152: out<=1;
   34153: out<=0;
   34154: out<=1;
   34155: out<=0;
   34156: out<=1;
   34157: out<=1;
   34158: out<=0;
   34159: out<=0;
   34160: out<=0;
   34161: out<=0;
   34162: out<=0;
   34163: out<=0;
   34164: out<=0;
   34165: out<=1;
   34166: out<=1;
   34167: out<=0;
   34168: out<=1;
   34169: out<=0;
   34170: out<=1;
   34171: out<=0;
   34172: out<=1;
   34173: out<=1;
   34174: out<=0;
   34175: out<=0;
   34176: out<=1;
   34177: out<=1;
   34178: out<=1;
   34179: out<=1;
   34180: out<=1;
   34181: out<=0;
   34182: out<=0;
   34183: out<=1;
   34184: out<=0;
   34185: out<=1;
   34186: out<=0;
   34187: out<=1;
   34188: out<=0;
   34189: out<=0;
   34190: out<=1;
   34191: out<=1;
   34192: out<=1;
   34193: out<=1;
   34194: out<=1;
   34195: out<=1;
   34196: out<=1;
   34197: out<=0;
   34198: out<=0;
   34199: out<=1;
   34200: out<=0;
   34201: out<=1;
   34202: out<=0;
   34203: out<=1;
   34204: out<=0;
   34205: out<=0;
   34206: out<=1;
   34207: out<=1;
   34208: out<=0;
   34209: out<=0;
   34210: out<=0;
   34211: out<=0;
   34212: out<=0;
   34213: out<=1;
   34214: out<=1;
   34215: out<=0;
   34216: out<=1;
   34217: out<=0;
   34218: out<=1;
   34219: out<=0;
   34220: out<=1;
   34221: out<=1;
   34222: out<=0;
   34223: out<=0;
   34224: out<=0;
   34225: out<=0;
   34226: out<=0;
   34227: out<=0;
   34228: out<=0;
   34229: out<=1;
   34230: out<=1;
   34231: out<=0;
   34232: out<=1;
   34233: out<=0;
   34234: out<=1;
   34235: out<=0;
   34236: out<=1;
   34237: out<=1;
   34238: out<=0;
   34239: out<=0;
   34240: out<=0;
   34241: out<=0;
   34242: out<=0;
   34243: out<=0;
   34244: out<=0;
   34245: out<=1;
   34246: out<=1;
   34247: out<=0;
   34248: out<=1;
   34249: out<=0;
   34250: out<=1;
   34251: out<=0;
   34252: out<=1;
   34253: out<=1;
   34254: out<=0;
   34255: out<=0;
   34256: out<=1;
   34257: out<=1;
   34258: out<=1;
   34259: out<=1;
   34260: out<=1;
   34261: out<=0;
   34262: out<=0;
   34263: out<=1;
   34264: out<=0;
   34265: out<=1;
   34266: out<=0;
   34267: out<=1;
   34268: out<=0;
   34269: out<=0;
   34270: out<=1;
   34271: out<=1;
   34272: out<=0;
   34273: out<=0;
   34274: out<=0;
   34275: out<=0;
   34276: out<=0;
   34277: out<=1;
   34278: out<=1;
   34279: out<=0;
   34280: out<=1;
   34281: out<=0;
   34282: out<=1;
   34283: out<=0;
   34284: out<=1;
   34285: out<=1;
   34286: out<=0;
   34287: out<=0;
   34288: out<=1;
   34289: out<=1;
   34290: out<=1;
   34291: out<=1;
   34292: out<=1;
   34293: out<=0;
   34294: out<=0;
   34295: out<=1;
   34296: out<=0;
   34297: out<=1;
   34298: out<=0;
   34299: out<=1;
   34300: out<=0;
   34301: out<=0;
   34302: out<=1;
   34303: out<=1;
   34304: out<=1;
   34305: out<=1;
   34306: out<=0;
   34307: out<=0;
   34308: out<=1;
   34309: out<=0;
   34310: out<=1;
   34311: out<=0;
   34312: out<=1;
   34313: out<=0;
   34314: out<=0;
   34315: out<=1;
   34316: out<=1;
   34317: out<=1;
   34318: out<=1;
   34319: out<=1;
   34320: out<=0;
   34321: out<=0;
   34322: out<=1;
   34323: out<=1;
   34324: out<=0;
   34325: out<=1;
   34326: out<=0;
   34327: out<=1;
   34328: out<=0;
   34329: out<=1;
   34330: out<=1;
   34331: out<=0;
   34332: out<=0;
   34333: out<=0;
   34334: out<=0;
   34335: out<=0;
   34336: out<=1;
   34337: out<=1;
   34338: out<=0;
   34339: out<=0;
   34340: out<=1;
   34341: out<=0;
   34342: out<=1;
   34343: out<=0;
   34344: out<=1;
   34345: out<=0;
   34346: out<=0;
   34347: out<=1;
   34348: out<=1;
   34349: out<=1;
   34350: out<=1;
   34351: out<=1;
   34352: out<=0;
   34353: out<=0;
   34354: out<=1;
   34355: out<=1;
   34356: out<=0;
   34357: out<=1;
   34358: out<=0;
   34359: out<=1;
   34360: out<=0;
   34361: out<=1;
   34362: out<=1;
   34363: out<=0;
   34364: out<=0;
   34365: out<=0;
   34366: out<=0;
   34367: out<=0;
   34368: out<=0;
   34369: out<=0;
   34370: out<=1;
   34371: out<=1;
   34372: out<=0;
   34373: out<=1;
   34374: out<=0;
   34375: out<=1;
   34376: out<=0;
   34377: out<=1;
   34378: out<=1;
   34379: out<=0;
   34380: out<=0;
   34381: out<=0;
   34382: out<=0;
   34383: out<=0;
   34384: out<=0;
   34385: out<=0;
   34386: out<=1;
   34387: out<=1;
   34388: out<=0;
   34389: out<=1;
   34390: out<=0;
   34391: out<=1;
   34392: out<=0;
   34393: out<=1;
   34394: out<=1;
   34395: out<=0;
   34396: out<=0;
   34397: out<=0;
   34398: out<=0;
   34399: out<=0;
   34400: out<=1;
   34401: out<=1;
   34402: out<=0;
   34403: out<=0;
   34404: out<=1;
   34405: out<=0;
   34406: out<=1;
   34407: out<=0;
   34408: out<=1;
   34409: out<=0;
   34410: out<=0;
   34411: out<=1;
   34412: out<=1;
   34413: out<=1;
   34414: out<=1;
   34415: out<=1;
   34416: out<=1;
   34417: out<=1;
   34418: out<=0;
   34419: out<=0;
   34420: out<=1;
   34421: out<=0;
   34422: out<=1;
   34423: out<=0;
   34424: out<=1;
   34425: out<=0;
   34426: out<=0;
   34427: out<=1;
   34428: out<=1;
   34429: out<=1;
   34430: out<=1;
   34431: out<=1;
   34432: out<=1;
   34433: out<=1;
   34434: out<=0;
   34435: out<=0;
   34436: out<=1;
   34437: out<=0;
   34438: out<=1;
   34439: out<=0;
   34440: out<=1;
   34441: out<=0;
   34442: out<=0;
   34443: out<=1;
   34444: out<=1;
   34445: out<=1;
   34446: out<=1;
   34447: out<=1;
   34448: out<=1;
   34449: out<=1;
   34450: out<=0;
   34451: out<=0;
   34452: out<=1;
   34453: out<=0;
   34454: out<=1;
   34455: out<=0;
   34456: out<=1;
   34457: out<=0;
   34458: out<=0;
   34459: out<=1;
   34460: out<=1;
   34461: out<=1;
   34462: out<=1;
   34463: out<=1;
   34464: out<=1;
   34465: out<=1;
   34466: out<=0;
   34467: out<=0;
   34468: out<=1;
   34469: out<=0;
   34470: out<=1;
   34471: out<=0;
   34472: out<=1;
   34473: out<=0;
   34474: out<=0;
   34475: out<=1;
   34476: out<=1;
   34477: out<=1;
   34478: out<=1;
   34479: out<=1;
   34480: out<=1;
   34481: out<=1;
   34482: out<=0;
   34483: out<=0;
   34484: out<=1;
   34485: out<=0;
   34486: out<=1;
   34487: out<=0;
   34488: out<=1;
   34489: out<=0;
   34490: out<=0;
   34491: out<=1;
   34492: out<=1;
   34493: out<=1;
   34494: out<=1;
   34495: out<=1;
   34496: out<=0;
   34497: out<=0;
   34498: out<=1;
   34499: out<=1;
   34500: out<=0;
   34501: out<=1;
   34502: out<=0;
   34503: out<=1;
   34504: out<=0;
   34505: out<=1;
   34506: out<=1;
   34507: out<=0;
   34508: out<=0;
   34509: out<=0;
   34510: out<=0;
   34511: out<=0;
   34512: out<=1;
   34513: out<=1;
   34514: out<=0;
   34515: out<=0;
   34516: out<=1;
   34517: out<=0;
   34518: out<=1;
   34519: out<=0;
   34520: out<=1;
   34521: out<=0;
   34522: out<=0;
   34523: out<=1;
   34524: out<=1;
   34525: out<=1;
   34526: out<=1;
   34527: out<=1;
   34528: out<=1;
   34529: out<=1;
   34530: out<=0;
   34531: out<=0;
   34532: out<=1;
   34533: out<=0;
   34534: out<=1;
   34535: out<=0;
   34536: out<=1;
   34537: out<=0;
   34538: out<=0;
   34539: out<=1;
   34540: out<=1;
   34541: out<=1;
   34542: out<=1;
   34543: out<=1;
   34544: out<=0;
   34545: out<=0;
   34546: out<=1;
   34547: out<=1;
   34548: out<=0;
   34549: out<=1;
   34550: out<=0;
   34551: out<=1;
   34552: out<=0;
   34553: out<=1;
   34554: out<=1;
   34555: out<=0;
   34556: out<=0;
   34557: out<=0;
   34558: out<=0;
   34559: out<=0;
   34560: out<=0;
   34561: out<=1;
   34562: out<=0;
   34563: out<=1;
   34564: out<=1;
   34565: out<=1;
   34566: out<=0;
   34567: out<=0;
   34568: out<=1;
   34569: out<=1;
   34570: out<=1;
   34571: out<=1;
   34572: out<=0;
   34573: out<=1;
   34574: out<=1;
   34575: out<=0;
   34576: out<=0;
   34577: out<=1;
   34578: out<=0;
   34579: out<=1;
   34580: out<=1;
   34581: out<=1;
   34582: out<=0;
   34583: out<=0;
   34584: out<=1;
   34585: out<=1;
   34586: out<=1;
   34587: out<=1;
   34588: out<=0;
   34589: out<=1;
   34590: out<=1;
   34591: out<=0;
   34592: out<=1;
   34593: out<=0;
   34594: out<=1;
   34595: out<=0;
   34596: out<=0;
   34597: out<=0;
   34598: out<=1;
   34599: out<=1;
   34600: out<=0;
   34601: out<=0;
   34602: out<=0;
   34603: out<=0;
   34604: out<=1;
   34605: out<=0;
   34606: out<=0;
   34607: out<=1;
   34608: out<=1;
   34609: out<=0;
   34610: out<=1;
   34611: out<=0;
   34612: out<=0;
   34613: out<=0;
   34614: out<=1;
   34615: out<=1;
   34616: out<=0;
   34617: out<=0;
   34618: out<=0;
   34619: out<=0;
   34620: out<=1;
   34621: out<=0;
   34622: out<=0;
   34623: out<=1;
   34624: out<=1;
   34625: out<=0;
   34626: out<=1;
   34627: out<=0;
   34628: out<=0;
   34629: out<=0;
   34630: out<=1;
   34631: out<=1;
   34632: out<=0;
   34633: out<=0;
   34634: out<=0;
   34635: out<=0;
   34636: out<=1;
   34637: out<=0;
   34638: out<=0;
   34639: out<=1;
   34640: out<=0;
   34641: out<=1;
   34642: out<=0;
   34643: out<=1;
   34644: out<=1;
   34645: out<=1;
   34646: out<=0;
   34647: out<=0;
   34648: out<=1;
   34649: out<=1;
   34650: out<=1;
   34651: out<=1;
   34652: out<=0;
   34653: out<=1;
   34654: out<=1;
   34655: out<=0;
   34656: out<=1;
   34657: out<=0;
   34658: out<=1;
   34659: out<=0;
   34660: out<=0;
   34661: out<=0;
   34662: out<=1;
   34663: out<=1;
   34664: out<=0;
   34665: out<=0;
   34666: out<=0;
   34667: out<=0;
   34668: out<=1;
   34669: out<=0;
   34670: out<=0;
   34671: out<=1;
   34672: out<=0;
   34673: out<=1;
   34674: out<=0;
   34675: out<=1;
   34676: out<=1;
   34677: out<=1;
   34678: out<=0;
   34679: out<=0;
   34680: out<=1;
   34681: out<=1;
   34682: out<=1;
   34683: out<=1;
   34684: out<=0;
   34685: out<=1;
   34686: out<=1;
   34687: out<=0;
   34688: out<=0;
   34689: out<=1;
   34690: out<=0;
   34691: out<=1;
   34692: out<=1;
   34693: out<=1;
   34694: out<=0;
   34695: out<=0;
   34696: out<=1;
   34697: out<=1;
   34698: out<=1;
   34699: out<=1;
   34700: out<=0;
   34701: out<=1;
   34702: out<=1;
   34703: out<=0;
   34704: out<=1;
   34705: out<=0;
   34706: out<=1;
   34707: out<=0;
   34708: out<=0;
   34709: out<=0;
   34710: out<=1;
   34711: out<=1;
   34712: out<=0;
   34713: out<=0;
   34714: out<=0;
   34715: out<=0;
   34716: out<=1;
   34717: out<=0;
   34718: out<=0;
   34719: out<=1;
   34720: out<=1;
   34721: out<=0;
   34722: out<=1;
   34723: out<=0;
   34724: out<=0;
   34725: out<=0;
   34726: out<=1;
   34727: out<=1;
   34728: out<=0;
   34729: out<=0;
   34730: out<=0;
   34731: out<=0;
   34732: out<=1;
   34733: out<=0;
   34734: out<=0;
   34735: out<=1;
   34736: out<=0;
   34737: out<=1;
   34738: out<=0;
   34739: out<=1;
   34740: out<=1;
   34741: out<=1;
   34742: out<=0;
   34743: out<=0;
   34744: out<=1;
   34745: out<=1;
   34746: out<=1;
   34747: out<=1;
   34748: out<=0;
   34749: out<=1;
   34750: out<=1;
   34751: out<=0;
   34752: out<=1;
   34753: out<=0;
   34754: out<=1;
   34755: out<=0;
   34756: out<=0;
   34757: out<=0;
   34758: out<=1;
   34759: out<=1;
   34760: out<=0;
   34761: out<=0;
   34762: out<=0;
   34763: out<=0;
   34764: out<=1;
   34765: out<=0;
   34766: out<=0;
   34767: out<=1;
   34768: out<=1;
   34769: out<=0;
   34770: out<=1;
   34771: out<=0;
   34772: out<=0;
   34773: out<=0;
   34774: out<=1;
   34775: out<=1;
   34776: out<=0;
   34777: out<=0;
   34778: out<=0;
   34779: out<=0;
   34780: out<=1;
   34781: out<=0;
   34782: out<=0;
   34783: out<=1;
   34784: out<=1;
   34785: out<=0;
   34786: out<=1;
   34787: out<=0;
   34788: out<=0;
   34789: out<=0;
   34790: out<=1;
   34791: out<=1;
   34792: out<=0;
   34793: out<=0;
   34794: out<=0;
   34795: out<=0;
   34796: out<=1;
   34797: out<=0;
   34798: out<=0;
   34799: out<=1;
   34800: out<=1;
   34801: out<=0;
   34802: out<=1;
   34803: out<=0;
   34804: out<=0;
   34805: out<=0;
   34806: out<=1;
   34807: out<=1;
   34808: out<=0;
   34809: out<=0;
   34810: out<=0;
   34811: out<=0;
   34812: out<=1;
   34813: out<=0;
   34814: out<=0;
   34815: out<=1;
   34816: out<=0;
   34817: out<=1;
   34818: out<=0;
   34819: out<=1;
   34820: out<=1;
   34821: out<=1;
   34822: out<=0;
   34823: out<=0;
   34824: out<=0;
   34825: out<=0;
   34826: out<=0;
   34827: out<=0;
   34828: out<=1;
   34829: out<=0;
   34830: out<=0;
   34831: out<=1;
   34832: out<=0;
   34833: out<=1;
   34834: out<=0;
   34835: out<=1;
   34836: out<=1;
   34837: out<=1;
   34838: out<=0;
   34839: out<=0;
   34840: out<=0;
   34841: out<=0;
   34842: out<=0;
   34843: out<=0;
   34844: out<=1;
   34845: out<=0;
   34846: out<=0;
   34847: out<=1;
   34848: out<=0;
   34849: out<=1;
   34850: out<=0;
   34851: out<=1;
   34852: out<=1;
   34853: out<=1;
   34854: out<=0;
   34855: out<=0;
   34856: out<=0;
   34857: out<=0;
   34858: out<=0;
   34859: out<=0;
   34860: out<=1;
   34861: out<=0;
   34862: out<=0;
   34863: out<=1;
   34864: out<=0;
   34865: out<=1;
   34866: out<=0;
   34867: out<=1;
   34868: out<=1;
   34869: out<=1;
   34870: out<=0;
   34871: out<=0;
   34872: out<=0;
   34873: out<=0;
   34874: out<=0;
   34875: out<=0;
   34876: out<=1;
   34877: out<=0;
   34878: out<=0;
   34879: out<=1;
   34880: out<=1;
   34881: out<=0;
   34882: out<=1;
   34883: out<=0;
   34884: out<=0;
   34885: out<=0;
   34886: out<=1;
   34887: out<=1;
   34888: out<=1;
   34889: out<=1;
   34890: out<=1;
   34891: out<=1;
   34892: out<=0;
   34893: out<=1;
   34894: out<=1;
   34895: out<=0;
   34896: out<=0;
   34897: out<=1;
   34898: out<=0;
   34899: out<=1;
   34900: out<=1;
   34901: out<=1;
   34902: out<=0;
   34903: out<=0;
   34904: out<=0;
   34905: out<=0;
   34906: out<=0;
   34907: out<=0;
   34908: out<=1;
   34909: out<=0;
   34910: out<=0;
   34911: out<=1;
   34912: out<=0;
   34913: out<=1;
   34914: out<=0;
   34915: out<=1;
   34916: out<=1;
   34917: out<=1;
   34918: out<=0;
   34919: out<=0;
   34920: out<=0;
   34921: out<=0;
   34922: out<=0;
   34923: out<=0;
   34924: out<=1;
   34925: out<=0;
   34926: out<=0;
   34927: out<=1;
   34928: out<=1;
   34929: out<=0;
   34930: out<=1;
   34931: out<=0;
   34932: out<=0;
   34933: out<=0;
   34934: out<=1;
   34935: out<=1;
   34936: out<=1;
   34937: out<=1;
   34938: out<=1;
   34939: out<=1;
   34940: out<=0;
   34941: out<=1;
   34942: out<=1;
   34943: out<=0;
   34944: out<=0;
   34945: out<=1;
   34946: out<=0;
   34947: out<=1;
   34948: out<=1;
   34949: out<=1;
   34950: out<=0;
   34951: out<=0;
   34952: out<=0;
   34953: out<=0;
   34954: out<=0;
   34955: out<=0;
   34956: out<=1;
   34957: out<=0;
   34958: out<=0;
   34959: out<=1;
   34960: out<=1;
   34961: out<=0;
   34962: out<=1;
   34963: out<=0;
   34964: out<=0;
   34965: out<=0;
   34966: out<=1;
   34967: out<=1;
   34968: out<=1;
   34969: out<=1;
   34970: out<=1;
   34971: out<=1;
   34972: out<=0;
   34973: out<=1;
   34974: out<=1;
   34975: out<=0;
   34976: out<=0;
   34977: out<=1;
   34978: out<=0;
   34979: out<=1;
   34980: out<=1;
   34981: out<=1;
   34982: out<=0;
   34983: out<=0;
   34984: out<=0;
   34985: out<=0;
   34986: out<=0;
   34987: out<=0;
   34988: out<=1;
   34989: out<=0;
   34990: out<=0;
   34991: out<=1;
   34992: out<=1;
   34993: out<=0;
   34994: out<=1;
   34995: out<=0;
   34996: out<=0;
   34997: out<=0;
   34998: out<=1;
   34999: out<=1;
   35000: out<=1;
   35001: out<=1;
   35002: out<=1;
   35003: out<=1;
   35004: out<=0;
   35005: out<=1;
   35006: out<=1;
   35007: out<=0;
   35008: out<=1;
   35009: out<=0;
   35010: out<=1;
   35011: out<=0;
   35012: out<=0;
   35013: out<=0;
   35014: out<=1;
   35015: out<=1;
   35016: out<=1;
   35017: out<=1;
   35018: out<=1;
   35019: out<=1;
   35020: out<=0;
   35021: out<=1;
   35022: out<=1;
   35023: out<=0;
   35024: out<=1;
   35025: out<=0;
   35026: out<=1;
   35027: out<=0;
   35028: out<=0;
   35029: out<=0;
   35030: out<=1;
   35031: out<=1;
   35032: out<=1;
   35033: out<=1;
   35034: out<=1;
   35035: out<=1;
   35036: out<=0;
   35037: out<=1;
   35038: out<=1;
   35039: out<=0;
   35040: out<=0;
   35041: out<=1;
   35042: out<=0;
   35043: out<=1;
   35044: out<=1;
   35045: out<=1;
   35046: out<=0;
   35047: out<=0;
   35048: out<=0;
   35049: out<=0;
   35050: out<=0;
   35051: out<=0;
   35052: out<=1;
   35053: out<=0;
   35054: out<=0;
   35055: out<=1;
   35056: out<=0;
   35057: out<=1;
   35058: out<=0;
   35059: out<=1;
   35060: out<=1;
   35061: out<=1;
   35062: out<=0;
   35063: out<=0;
   35064: out<=0;
   35065: out<=0;
   35066: out<=0;
   35067: out<=0;
   35068: out<=1;
   35069: out<=0;
   35070: out<=0;
   35071: out<=1;
   35072: out<=1;
   35073: out<=1;
   35074: out<=0;
   35075: out<=0;
   35076: out<=1;
   35077: out<=0;
   35078: out<=1;
   35079: out<=0;
   35080: out<=0;
   35081: out<=1;
   35082: out<=1;
   35083: out<=0;
   35084: out<=0;
   35085: out<=0;
   35086: out<=0;
   35087: out<=0;
   35088: out<=0;
   35089: out<=0;
   35090: out<=1;
   35091: out<=1;
   35092: out<=0;
   35093: out<=1;
   35094: out<=0;
   35095: out<=1;
   35096: out<=1;
   35097: out<=0;
   35098: out<=0;
   35099: out<=1;
   35100: out<=1;
   35101: out<=1;
   35102: out<=1;
   35103: out<=1;
   35104: out<=0;
   35105: out<=0;
   35106: out<=1;
   35107: out<=1;
   35108: out<=0;
   35109: out<=1;
   35110: out<=0;
   35111: out<=1;
   35112: out<=1;
   35113: out<=0;
   35114: out<=0;
   35115: out<=1;
   35116: out<=1;
   35117: out<=1;
   35118: out<=1;
   35119: out<=1;
   35120: out<=1;
   35121: out<=1;
   35122: out<=0;
   35123: out<=0;
   35124: out<=1;
   35125: out<=0;
   35126: out<=1;
   35127: out<=0;
   35128: out<=0;
   35129: out<=1;
   35130: out<=1;
   35131: out<=0;
   35132: out<=0;
   35133: out<=0;
   35134: out<=0;
   35135: out<=0;
   35136: out<=0;
   35137: out<=0;
   35138: out<=1;
   35139: out<=1;
   35140: out<=0;
   35141: out<=1;
   35142: out<=0;
   35143: out<=1;
   35144: out<=1;
   35145: out<=0;
   35146: out<=0;
   35147: out<=1;
   35148: out<=1;
   35149: out<=1;
   35150: out<=1;
   35151: out<=1;
   35152: out<=0;
   35153: out<=0;
   35154: out<=1;
   35155: out<=1;
   35156: out<=0;
   35157: out<=1;
   35158: out<=0;
   35159: out<=1;
   35160: out<=1;
   35161: out<=0;
   35162: out<=0;
   35163: out<=1;
   35164: out<=1;
   35165: out<=1;
   35166: out<=1;
   35167: out<=1;
   35168: out<=0;
   35169: out<=0;
   35170: out<=1;
   35171: out<=1;
   35172: out<=0;
   35173: out<=1;
   35174: out<=0;
   35175: out<=1;
   35176: out<=1;
   35177: out<=0;
   35178: out<=0;
   35179: out<=1;
   35180: out<=1;
   35181: out<=1;
   35182: out<=1;
   35183: out<=1;
   35184: out<=0;
   35185: out<=0;
   35186: out<=1;
   35187: out<=1;
   35188: out<=0;
   35189: out<=1;
   35190: out<=0;
   35191: out<=1;
   35192: out<=1;
   35193: out<=0;
   35194: out<=0;
   35195: out<=1;
   35196: out<=1;
   35197: out<=1;
   35198: out<=1;
   35199: out<=1;
   35200: out<=1;
   35201: out<=1;
   35202: out<=0;
   35203: out<=0;
   35204: out<=1;
   35205: out<=0;
   35206: out<=1;
   35207: out<=0;
   35208: out<=0;
   35209: out<=1;
   35210: out<=1;
   35211: out<=0;
   35212: out<=0;
   35213: out<=0;
   35214: out<=0;
   35215: out<=0;
   35216: out<=1;
   35217: out<=1;
   35218: out<=0;
   35219: out<=0;
   35220: out<=1;
   35221: out<=0;
   35222: out<=1;
   35223: out<=0;
   35224: out<=0;
   35225: out<=1;
   35226: out<=1;
   35227: out<=0;
   35228: out<=0;
   35229: out<=0;
   35230: out<=0;
   35231: out<=0;
   35232: out<=0;
   35233: out<=0;
   35234: out<=1;
   35235: out<=1;
   35236: out<=0;
   35237: out<=1;
   35238: out<=0;
   35239: out<=1;
   35240: out<=1;
   35241: out<=0;
   35242: out<=0;
   35243: out<=1;
   35244: out<=1;
   35245: out<=1;
   35246: out<=1;
   35247: out<=1;
   35248: out<=0;
   35249: out<=0;
   35250: out<=1;
   35251: out<=1;
   35252: out<=0;
   35253: out<=1;
   35254: out<=0;
   35255: out<=1;
   35256: out<=1;
   35257: out<=0;
   35258: out<=0;
   35259: out<=1;
   35260: out<=1;
   35261: out<=1;
   35262: out<=1;
   35263: out<=1;
   35264: out<=0;
   35265: out<=0;
   35266: out<=1;
   35267: out<=1;
   35268: out<=0;
   35269: out<=1;
   35270: out<=0;
   35271: out<=1;
   35272: out<=1;
   35273: out<=0;
   35274: out<=0;
   35275: out<=1;
   35276: out<=1;
   35277: out<=1;
   35278: out<=1;
   35279: out<=1;
   35280: out<=1;
   35281: out<=1;
   35282: out<=0;
   35283: out<=0;
   35284: out<=1;
   35285: out<=0;
   35286: out<=1;
   35287: out<=0;
   35288: out<=0;
   35289: out<=1;
   35290: out<=1;
   35291: out<=0;
   35292: out<=0;
   35293: out<=0;
   35294: out<=0;
   35295: out<=0;
   35296: out<=0;
   35297: out<=0;
   35298: out<=1;
   35299: out<=1;
   35300: out<=0;
   35301: out<=1;
   35302: out<=0;
   35303: out<=1;
   35304: out<=1;
   35305: out<=0;
   35306: out<=0;
   35307: out<=1;
   35308: out<=1;
   35309: out<=1;
   35310: out<=1;
   35311: out<=1;
   35312: out<=1;
   35313: out<=1;
   35314: out<=0;
   35315: out<=0;
   35316: out<=1;
   35317: out<=0;
   35318: out<=1;
   35319: out<=0;
   35320: out<=0;
   35321: out<=1;
   35322: out<=1;
   35323: out<=0;
   35324: out<=0;
   35325: out<=0;
   35326: out<=0;
   35327: out<=0;
   35328: out<=0;
   35329: out<=0;
   35330: out<=0;
   35331: out<=0;
   35332: out<=0;
   35333: out<=1;
   35334: out<=1;
   35335: out<=0;
   35336: out<=0;
   35337: out<=1;
   35338: out<=0;
   35339: out<=1;
   35340: out<=0;
   35341: out<=0;
   35342: out<=1;
   35343: out<=1;
   35344: out<=1;
   35345: out<=1;
   35346: out<=1;
   35347: out<=1;
   35348: out<=1;
   35349: out<=0;
   35350: out<=0;
   35351: out<=1;
   35352: out<=1;
   35353: out<=0;
   35354: out<=1;
   35355: out<=0;
   35356: out<=1;
   35357: out<=1;
   35358: out<=0;
   35359: out<=0;
   35360: out<=0;
   35361: out<=0;
   35362: out<=0;
   35363: out<=0;
   35364: out<=0;
   35365: out<=1;
   35366: out<=1;
   35367: out<=0;
   35368: out<=0;
   35369: out<=1;
   35370: out<=0;
   35371: out<=1;
   35372: out<=0;
   35373: out<=0;
   35374: out<=1;
   35375: out<=1;
   35376: out<=1;
   35377: out<=1;
   35378: out<=1;
   35379: out<=1;
   35380: out<=1;
   35381: out<=0;
   35382: out<=0;
   35383: out<=1;
   35384: out<=1;
   35385: out<=0;
   35386: out<=1;
   35387: out<=0;
   35388: out<=1;
   35389: out<=1;
   35390: out<=0;
   35391: out<=0;
   35392: out<=1;
   35393: out<=1;
   35394: out<=1;
   35395: out<=1;
   35396: out<=1;
   35397: out<=0;
   35398: out<=0;
   35399: out<=1;
   35400: out<=1;
   35401: out<=0;
   35402: out<=1;
   35403: out<=0;
   35404: out<=1;
   35405: out<=1;
   35406: out<=0;
   35407: out<=0;
   35408: out<=1;
   35409: out<=1;
   35410: out<=1;
   35411: out<=1;
   35412: out<=1;
   35413: out<=0;
   35414: out<=0;
   35415: out<=1;
   35416: out<=1;
   35417: out<=0;
   35418: out<=1;
   35419: out<=0;
   35420: out<=1;
   35421: out<=1;
   35422: out<=0;
   35423: out<=0;
   35424: out<=0;
   35425: out<=0;
   35426: out<=0;
   35427: out<=0;
   35428: out<=0;
   35429: out<=1;
   35430: out<=1;
   35431: out<=0;
   35432: out<=0;
   35433: out<=1;
   35434: out<=0;
   35435: out<=1;
   35436: out<=0;
   35437: out<=0;
   35438: out<=1;
   35439: out<=1;
   35440: out<=0;
   35441: out<=0;
   35442: out<=0;
   35443: out<=0;
   35444: out<=0;
   35445: out<=1;
   35446: out<=1;
   35447: out<=0;
   35448: out<=0;
   35449: out<=1;
   35450: out<=0;
   35451: out<=1;
   35452: out<=0;
   35453: out<=0;
   35454: out<=1;
   35455: out<=1;
   35456: out<=0;
   35457: out<=0;
   35458: out<=0;
   35459: out<=0;
   35460: out<=0;
   35461: out<=1;
   35462: out<=1;
   35463: out<=0;
   35464: out<=0;
   35465: out<=1;
   35466: out<=0;
   35467: out<=1;
   35468: out<=0;
   35469: out<=0;
   35470: out<=1;
   35471: out<=1;
   35472: out<=0;
   35473: out<=0;
   35474: out<=0;
   35475: out<=0;
   35476: out<=0;
   35477: out<=1;
   35478: out<=1;
   35479: out<=0;
   35480: out<=0;
   35481: out<=1;
   35482: out<=0;
   35483: out<=1;
   35484: out<=0;
   35485: out<=0;
   35486: out<=1;
   35487: out<=1;
   35488: out<=0;
   35489: out<=0;
   35490: out<=0;
   35491: out<=0;
   35492: out<=0;
   35493: out<=1;
   35494: out<=1;
   35495: out<=0;
   35496: out<=0;
   35497: out<=1;
   35498: out<=0;
   35499: out<=1;
   35500: out<=0;
   35501: out<=0;
   35502: out<=1;
   35503: out<=1;
   35504: out<=0;
   35505: out<=0;
   35506: out<=0;
   35507: out<=0;
   35508: out<=0;
   35509: out<=1;
   35510: out<=1;
   35511: out<=0;
   35512: out<=0;
   35513: out<=1;
   35514: out<=0;
   35515: out<=1;
   35516: out<=0;
   35517: out<=0;
   35518: out<=1;
   35519: out<=1;
   35520: out<=1;
   35521: out<=1;
   35522: out<=1;
   35523: out<=1;
   35524: out<=1;
   35525: out<=0;
   35526: out<=0;
   35527: out<=1;
   35528: out<=1;
   35529: out<=0;
   35530: out<=1;
   35531: out<=0;
   35532: out<=1;
   35533: out<=1;
   35534: out<=0;
   35535: out<=0;
   35536: out<=0;
   35537: out<=0;
   35538: out<=0;
   35539: out<=0;
   35540: out<=0;
   35541: out<=1;
   35542: out<=1;
   35543: out<=0;
   35544: out<=0;
   35545: out<=1;
   35546: out<=0;
   35547: out<=1;
   35548: out<=0;
   35549: out<=0;
   35550: out<=1;
   35551: out<=1;
   35552: out<=0;
   35553: out<=0;
   35554: out<=0;
   35555: out<=0;
   35556: out<=0;
   35557: out<=1;
   35558: out<=1;
   35559: out<=0;
   35560: out<=0;
   35561: out<=1;
   35562: out<=0;
   35563: out<=1;
   35564: out<=0;
   35565: out<=0;
   35566: out<=1;
   35567: out<=1;
   35568: out<=1;
   35569: out<=1;
   35570: out<=1;
   35571: out<=1;
   35572: out<=1;
   35573: out<=0;
   35574: out<=0;
   35575: out<=1;
   35576: out<=1;
   35577: out<=0;
   35578: out<=1;
   35579: out<=0;
   35580: out<=1;
   35581: out<=1;
   35582: out<=0;
   35583: out<=0;
   35584: out<=1;
   35585: out<=0;
   35586: out<=0;
   35587: out<=1;
   35588: out<=0;
   35589: out<=0;
   35590: out<=0;
   35591: out<=0;
   35592: out<=0;
   35593: out<=0;
   35594: out<=1;
   35595: out<=1;
   35596: out<=1;
   35597: out<=0;
   35598: out<=1;
   35599: out<=0;
   35600: out<=1;
   35601: out<=0;
   35602: out<=0;
   35603: out<=1;
   35604: out<=0;
   35605: out<=0;
   35606: out<=0;
   35607: out<=0;
   35608: out<=0;
   35609: out<=0;
   35610: out<=1;
   35611: out<=1;
   35612: out<=1;
   35613: out<=0;
   35614: out<=1;
   35615: out<=0;
   35616: out<=0;
   35617: out<=1;
   35618: out<=1;
   35619: out<=0;
   35620: out<=1;
   35621: out<=1;
   35622: out<=1;
   35623: out<=1;
   35624: out<=1;
   35625: out<=1;
   35626: out<=0;
   35627: out<=0;
   35628: out<=0;
   35629: out<=1;
   35630: out<=0;
   35631: out<=1;
   35632: out<=0;
   35633: out<=1;
   35634: out<=1;
   35635: out<=0;
   35636: out<=1;
   35637: out<=1;
   35638: out<=1;
   35639: out<=1;
   35640: out<=1;
   35641: out<=1;
   35642: out<=0;
   35643: out<=0;
   35644: out<=0;
   35645: out<=1;
   35646: out<=0;
   35647: out<=1;
   35648: out<=0;
   35649: out<=1;
   35650: out<=1;
   35651: out<=0;
   35652: out<=1;
   35653: out<=1;
   35654: out<=1;
   35655: out<=1;
   35656: out<=1;
   35657: out<=1;
   35658: out<=0;
   35659: out<=0;
   35660: out<=0;
   35661: out<=1;
   35662: out<=0;
   35663: out<=1;
   35664: out<=1;
   35665: out<=0;
   35666: out<=0;
   35667: out<=1;
   35668: out<=0;
   35669: out<=0;
   35670: out<=0;
   35671: out<=0;
   35672: out<=0;
   35673: out<=0;
   35674: out<=1;
   35675: out<=1;
   35676: out<=1;
   35677: out<=0;
   35678: out<=1;
   35679: out<=0;
   35680: out<=0;
   35681: out<=1;
   35682: out<=1;
   35683: out<=0;
   35684: out<=1;
   35685: out<=1;
   35686: out<=1;
   35687: out<=1;
   35688: out<=1;
   35689: out<=1;
   35690: out<=0;
   35691: out<=0;
   35692: out<=0;
   35693: out<=1;
   35694: out<=0;
   35695: out<=1;
   35696: out<=1;
   35697: out<=0;
   35698: out<=0;
   35699: out<=1;
   35700: out<=0;
   35701: out<=0;
   35702: out<=0;
   35703: out<=0;
   35704: out<=0;
   35705: out<=0;
   35706: out<=1;
   35707: out<=1;
   35708: out<=1;
   35709: out<=0;
   35710: out<=1;
   35711: out<=0;
   35712: out<=1;
   35713: out<=0;
   35714: out<=0;
   35715: out<=1;
   35716: out<=0;
   35717: out<=0;
   35718: out<=0;
   35719: out<=0;
   35720: out<=0;
   35721: out<=0;
   35722: out<=1;
   35723: out<=1;
   35724: out<=1;
   35725: out<=0;
   35726: out<=1;
   35727: out<=0;
   35728: out<=0;
   35729: out<=1;
   35730: out<=1;
   35731: out<=0;
   35732: out<=1;
   35733: out<=1;
   35734: out<=1;
   35735: out<=1;
   35736: out<=1;
   35737: out<=1;
   35738: out<=0;
   35739: out<=0;
   35740: out<=0;
   35741: out<=1;
   35742: out<=0;
   35743: out<=1;
   35744: out<=0;
   35745: out<=1;
   35746: out<=1;
   35747: out<=0;
   35748: out<=1;
   35749: out<=1;
   35750: out<=1;
   35751: out<=1;
   35752: out<=1;
   35753: out<=1;
   35754: out<=0;
   35755: out<=0;
   35756: out<=0;
   35757: out<=1;
   35758: out<=0;
   35759: out<=1;
   35760: out<=1;
   35761: out<=0;
   35762: out<=0;
   35763: out<=1;
   35764: out<=0;
   35765: out<=0;
   35766: out<=0;
   35767: out<=0;
   35768: out<=0;
   35769: out<=0;
   35770: out<=1;
   35771: out<=1;
   35772: out<=1;
   35773: out<=0;
   35774: out<=1;
   35775: out<=0;
   35776: out<=0;
   35777: out<=1;
   35778: out<=1;
   35779: out<=0;
   35780: out<=1;
   35781: out<=1;
   35782: out<=1;
   35783: out<=1;
   35784: out<=1;
   35785: out<=1;
   35786: out<=0;
   35787: out<=0;
   35788: out<=0;
   35789: out<=1;
   35790: out<=0;
   35791: out<=1;
   35792: out<=0;
   35793: out<=1;
   35794: out<=1;
   35795: out<=0;
   35796: out<=1;
   35797: out<=1;
   35798: out<=1;
   35799: out<=1;
   35800: out<=1;
   35801: out<=1;
   35802: out<=0;
   35803: out<=0;
   35804: out<=0;
   35805: out<=1;
   35806: out<=0;
   35807: out<=1;
   35808: out<=0;
   35809: out<=1;
   35810: out<=1;
   35811: out<=0;
   35812: out<=1;
   35813: out<=1;
   35814: out<=1;
   35815: out<=1;
   35816: out<=1;
   35817: out<=1;
   35818: out<=0;
   35819: out<=0;
   35820: out<=0;
   35821: out<=1;
   35822: out<=0;
   35823: out<=1;
   35824: out<=0;
   35825: out<=1;
   35826: out<=1;
   35827: out<=0;
   35828: out<=1;
   35829: out<=1;
   35830: out<=1;
   35831: out<=1;
   35832: out<=1;
   35833: out<=1;
   35834: out<=0;
   35835: out<=0;
   35836: out<=0;
   35837: out<=1;
   35838: out<=0;
   35839: out<=1;
   35840: out<=0;
   35841: out<=0;
   35842: out<=1;
   35843: out<=1;
   35844: out<=1;
   35845: out<=0;
   35846: out<=1;
   35847: out<=0;
   35848: out<=0;
   35849: out<=1;
   35850: out<=1;
   35851: out<=0;
   35852: out<=1;
   35853: out<=1;
   35854: out<=1;
   35855: out<=1;
   35856: out<=0;
   35857: out<=0;
   35858: out<=1;
   35859: out<=1;
   35860: out<=1;
   35861: out<=0;
   35862: out<=1;
   35863: out<=0;
   35864: out<=0;
   35865: out<=1;
   35866: out<=1;
   35867: out<=0;
   35868: out<=1;
   35869: out<=1;
   35870: out<=1;
   35871: out<=1;
   35872: out<=0;
   35873: out<=0;
   35874: out<=1;
   35875: out<=1;
   35876: out<=1;
   35877: out<=0;
   35878: out<=1;
   35879: out<=0;
   35880: out<=0;
   35881: out<=1;
   35882: out<=1;
   35883: out<=0;
   35884: out<=1;
   35885: out<=1;
   35886: out<=1;
   35887: out<=1;
   35888: out<=0;
   35889: out<=0;
   35890: out<=1;
   35891: out<=1;
   35892: out<=1;
   35893: out<=0;
   35894: out<=1;
   35895: out<=0;
   35896: out<=0;
   35897: out<=1;
   35898: out<=1;
   35899: out<=0;
   35900: out<=1;
   35901: out<=1;
   35902: out<=1;
   35903: out<=1;
   35904: out<=1;
   35905: out<=1;
   35906: out<=0;
   35907: out<=0;
   35908: out<=0;
   35909: out<=1;
   35910: out<=0;
   35911: out<=1;
   35912: out<=1;
   35913: out<=0;
   35914: out<=0;
   35915: out<=1;
   35916: out<=0;
   35917: out<=0;
   35918: out<=0;
   35919: out<=0;
   35920: out<=0;
   35921: out<=0;
   35922: out<=1;
   35923: out<=1;
   35924: out<=1;
   35925: out<=0;
   35926: out<=1;
   35927: out<=0;
   35928: out<=0;
   35929: out<=1;
   35930: out<=1;
   35931: out<=0;
   35932: out<=1;
   35933: out<=1;
   35934: out<=1;
   35935: out<=1;
   35936: out<=0;
   35937: out<=0;
   35938: out<=1;
   35939: out<=1;
   35940: out<=1;
   35941: out<=0;
   35942: out<=1;
   35943: out<=0;
   35944: out<=0;
   35945: out<=1;
   35946: out<=1;
   35947: out<=0;
   35948: out<=1;
   35949: out<=1;
   35950: out<=1;
   35951: out<=1;
   35952: out<=1;
   35953: out<=1;
   35954: out<=0;
   35955: out<=0;
   35956: out<=0;
   35957: out<=1;
   35958: out<=0;
   35959: out<=1;
   35960: out<=1;
   35961: out<=0;
   35962: out<=0;
   35963: out<=1;
   35964: out<=0;
   35965: out<=0;
   35966: out<=0;
   35967: out<=0;
   35968: out<=0;
   35969: out<=0;
   35970: out<=1;
   35971: out<=1;
   35972: out<=1;
   35973: out<=0;
   35974: out<=1;
   35975: out<=0;
   35976: out<=0;
   35977: out<=1;
   35978: out<=1;
   35979: out<=0;
   35980: out<=1;
   35981: out<=1;
   35982: out<=1;
   35983: out<=1;
   35984: out<=1;
   35985: out<=1;
   35986: out<=0;
   35987: out<=0;
   35988: out<=0;
   35989: out<=1;
   35990: out<=0;
   35991: out<=1;
   35992: out<=1;
   35993: out<=0;
   35994: out<=0;
   35995: out<=1;
   35996: out<=0;
   35997: out<=0;
   35998: out<=0;
   35999: out<=0;
   36000: out<=0;
   36001: out<=0;
   36002: out<=1;
   36003: out<=1;
   36004: out<=1;
   36005: out<=0;
   36006: out<=1;
   36007: out<=0;
   36008: out<=0;
   36009: out<=1;
   36010: out<=1;
   36011: out<=0;
   36012: out<=1;
   36013: out<=1;
   36014: out<=1;
   36015: out<=1;
   36016: out<=1;
   36017: out<=1;
   36018: out<=0;
   36019: out<=0;
   36020: out<=0;
   36021: out<=1;
   36022: out<=0;
   36023: out<=1;
   36024: out<=1;
   36025: out<=0;
   36026: out<=0;
   36027: out<=1;
   36028: out<=0;
   36029: out<=0;
   36030: out<=0;
   36031: out<=0;
   36032: out<=1;
   36033: out<=1;
   36034: out<=0;
   36035: out<=0;
   36036: out<=0;
   36037: out<=1;
   36038: out<=0;
   36039: out<=1;
   36040: out<=1;
   36041: out<=0;
   36042: out<=0;
   36043: out<=1;
   36044: out<=0;
   36045: out<=0;
   36046: out<=0;
   36047: out<=0;
   36048: out<=1;
   36049: out<=1;
   36050: out<=0;
   36051: out<=0;
   36052: out<=0;
   36053: out<=1;
   36054: out<=0;
   36055: out<=1;
   36056: out<=1;
   36057: out<=0;
   36058: out<=0;
   36059: out<=1;
   36060: out<=0;
   36061: out<=0;
   36062: out<=0;
   36063: out<=0;
   36064: out<=0;
   36065: out<=0;
   36066: out<=1;
   36067: out<=1;
   36068: out<=1;
   36069: out<=0;
   36070: out<=1;
   36071: out<=0;
   36072: out<=0;
   36073: out<=1;
   36074: out<=1;
   36075: out<=0;
   36076: out<=1;
   36077: out<=1;
   36078: out<=1;
   36079: out<=1;
   36080: out<=0;
   36081: out<=0;
   36082: out<=1;
   36083: out<=1;
   36084: out<=1;
   36085: out<=0;
   36086: out<=1;
   36087: out<=0;
   36088: out<=0;
   36089: out<=1;
   36090: out<=1;
   36091: out<=0;
   36092: out<=1;
   36093: out<=1;
   36094: out<=1;
   36095: out<=1;
   36096: out<=0;
   36097: out<=1;
   36098: out<=0;
   36099: out<=1;
   36100: out<=0;
   36101: out<=0;
   36102: out<=1;
   36103: out<=1;
   36104: out<=1;
   36105: out<=1;
   36106: out<=1;
   36107: out<=1;
   36108: out<=1;
   36109: out<=0;
   36110: out<=0;
   36111: out<=1;
   36112: out<=1;
   36113: out<=0;
   36114: out<=1;
   36115: out<=0;
   36116: out<=1;
   36117: out<=1;
   36118: out<=0;
   36119: out<=0;
   36120: out<=0;
   36121: out<=0;
   36122: out<=0;
   36123: out<=0;
   36124: out<=0;
   36125: out<=1;
   36126: out<=1;
   36127: out<=0;
   36128: out<=1;
   36129: out<=0;
   36130: out<=1;
   36131: out<=0;
   36132: out<=1;
   36133: out<=1;
   36134: out<=0;
   36135: out<=0;
   36136: out<=0;
   36137: out<=0;
   36138: out<=0;
   36139: out<=0;
   36140: out<=0;
   36141: out<=1;
   36142: out<=1;
   36143: out<=0;
   36144: out<=0;
   36145: out<=1;
   36146: out<=0;
   36147: out<=1;
   36148: out<=0;
   36149: out<=0;
   36150: out<=1;
   36151: out<=1;
   36152: out<=1;
   36153: out<=1;
   36154: out<=1;
   36155: out<=1;
   36156: out<=1;
   36157: out<=0;
   36158: out<=0;
   36159: out<=1;
   36160: out<=1;
   36161: out<=0;
   36162: out<=1;
   36163: out<=0;
   36164: out<=1;
   36165: out<=1;
   36166: out<=0;
   36167: out<=0;
   36168: out<=0;
   36169: out<=0;
   36170: out<=0;
   36171: out<=0;
   36172: out<=0;
   36173: out<=1;
   36174: out<=1;
   36175: out<=0;
   36176: out<=1;
   36177: out<=0;
   36178: out<=1;
   36179: out<=0;
   36180: out<=1;
   36181: out<=1;
   36182: out<=0;
   36183: out<=0;
   36184: out<=0;
   36185: out<=0;
   36186: out<=0;
   36187: out<=0;
   36188: out<=0;
   36189: out<=1;
   36190: out<=1;
   36191: out<=0;
   36192: out<=1;
   36193: out<=0;
   36194: out<=1;
   36195: out<=0;
   36196: out<=1;
   36197: out<=1;
   36198: out<=0;
   36199: out<=0;
   36200: out<=0;
   36201: out<=0;
   36202: out<=0;
   36203: out<=0;
   36204: out<=0;
   36205: out<=1;
   36206: out<=1;
   36207: out<=0;
   36208: out<=1;
   36209: out<=0;
   36210: out<=1;
   36211: out<=0;
   36212: out<=1;
   36213: out<=1;
   36214: out<=0;
   36215: out<=0;
   36216: out<=0;
   36217: out<=0;
   36218: out<=0;
   36219: out<=0;
   36220: out<=0;
   36221: out<=1;
   36222: out<=1;
   36223: out<=0;
   36224: out<=0;
   36225: out<=1;
   36226: out<=0;
   36227: out<=1;
   36228: out<=0;
   36229: out<=0;
   36230: out<=1;
   36231: out<=1;
   36232: out<=1;
   36233: out<=1;
   36234: out<=1;
   36235: out<=1;
   36236: out<=1;
   36237: out<=0;
   36238: out<=0;
   36239: out<=1;
   36240: out<=0;
   36241: out<=1;
   36242: out<=0;
   36243: out<=1;
   36244: out<=0;
   36245: out<=0;
   36246: out<=1;
   36247: out<=1;
   36248: out<=1;
   36249: out<=1;
   36250: out<=1;
   36251: out<=1;
   36252: out<=1;
   36253: out<=0;
   36254: out<=0;
   36255: out<=1;
   36256: out<=1;
   36257: out<=0;
   36258: out<=1;
   36259: out<=0;
   36260: out<=1;
   36261: out<=1;
   36262: out<=0;
   36263: out<=0;
   36264: out<=0;
   36265: out<=0;
   36266: out<=0;
   36267: out<=0;
   36268: out<=0;
   36269: out<=1;
   36270: out<=1;
   36271: out<=0;
   36272: out<=1;
   36273: out<=0;
   36274: out<=1;
   36275: out<=0;
   36276: out<=1;
   36277: out<=1;
   36278: out<=0;
   36279: out<=0;
   36280: out<=0;
   36281: out<=0;
   36282: out<=0;
   36283: out<=0;
   36284: out<=0;
   36285: out<=1;
   36286: out<=1;
   36287: out<=0;
   36288: out<=1;
   36289: out<=0;
   36290: out<=1;
   36291: out<=0;
   36292: out<=1;
   36293: out<=1;
   36294: out<=0;
   36295: out<=0;
   36296: out<=0;
   36297: out<=0;
   36298: out<=0;
   36299: out<=0;
   36300: out<=0;
   36301: out<=1;
   36302: out<=1;
   36303: out<=0;
   36304: out<=0;
   36305: out<=1;
   36306: out<=0;
   36307: out<=1;
   36308: out<=0;
   36309: out<=0;
   36310: out<=1;
   36311: out<=1;
   36312: out<=1;
   36313: out<=1;
   36314: out<=1;
   36315: out<=1;
   36316: out<=1;
   36317: out<=0;
   36318: out<=0;
   36319: out<=1;
   36320: out<=1;
   36321: out<=0;
   36322: out<=1;
   36323: out<=0;
   36324: out<=1;
   36325: out<=1;
   36326: out<=0;
   36327: out<=0;
   36328: out<=0;
   36329: out<=0;
   36330: out<=0;
   36331: out<=0;
   36332: out<=0;
   36333: out<=1;
   36334: out<=1;
   36335: out<=0;
   36336: out<=0;
   36337: out<=1;
   36338: out<=0;
   36339: out<=1;
   36340: out<=0;
   36341: out<=0;
   36342: out<=1;
   36343: out<=1;
   36344: out<=1;
   36345: out<=1;
   36346: out<=1;
   36347: out<=1;
   36348: out<=1;
   36349: out<=0;
   36350: out<=0;
   36351: out<=1;
   36352: out<=1;
   36353: out<=0;
   36354: out<=0;
   36355: out<=1;
   36356: out<=1;
   36357: out<=1;
   36358: out<=1;
   36359: out<=1;
   36360: out<=1;
   36361: out<=1;
   36362: out<=0;
   36363: out<=0;
   36364: out<=1;
   36365: out<=0;
   36366: out<=1;
   36367: out<=0;
   36368: out<=0;
   36369: out<=1;
   36370: out<=1;
   36371: out<=0;
   36372: out<=0;
   36373: out<=0;
   36374: out<=0;
   36375: out<=0;
   36376: out<=0;
   36377: out<=0;
   36378: out<=1;
   36379: out<=1;
   36380: out<=0;
   36381: out<=1;
   36382: out<=0;
   36383: out<=1;
   36384: out<=1;
   36385: out<=0;
   36386: out<=0;
   36387: out<=1;
   36388: out<=1;
   36389: out<=1;
   36390: out<=1;
   36391: out<=1;
   36392: out<=1;
   36393: out<=1;
   36394: out<=0;
   36395: out<=0;
   36396: out<=1;
   36397: out<=0;
   36398: out<=1;
   36399: out<=0;
   36400: out<=0;
   36401: out<=1;
   36402: out<=1;
   36403: out<=0;
   36404: out<=0;
   36405: out<=0;
   36406: out<=0;
   36407: out<=0;
   36408: out<=0;
   36409: out<=0;
   36410: out<=1;
   36411: out<=1;
   36412: out<=0;
   36413: out<=1;
   36414: out<=0;
   36415: out<=1;
   36416: out<=0;
   36417: out<=1;
   36418: out<=1;
   36419: out<=0;
   36420: out<=0;
   36421: out<=0;
   36422: out<=0;
   36423: out<=0;
   36424: out<=0;
   36425: out<=0;
   36426: out<=1;
   36427: out<=1;
   36428: out<=0;
   36429: out<=1;
   36430: out<=0;
   36431: out<=1;
   36432: out<=0;
   36433: out<=1;
   36434: out<=1;
   36435: out<=0;
   36436: out<=0;
   36437: out<=0;
   36438: out<=0;
   36439: out<=0;
   36440: out<=0;
   36441: out<=0;
   36442: out<=1;
   36443: out<=1;
   36444: out<=0;
   36445: out<=1;
   36446: out<=0;
   36447: out<=1;
   36448: out<=1;
   36449: out<=0;
   36450: out<=0;
   36451: out<=1;
   36452: out<=1;
   36453: out<=1;
   36454: out<=1;
   36455: out<=1;
   36456: out<=1;
   36457: out<=1;
   36458: out<=0;
   36459: out<=0;
   36460: out<=1;
   36461: out<=0;
   36462: out<=1;
   36463: out<=0;
   36464: out<=1;
   36465: out<=0;
   36466: out<=0;
   36467: out<=1;
   36468: out<=1;
   36469: out<=1;
   36470: out<=1;
   36471: out<=1;
   36472: out<=1;
   36473: out<=1;
   36474: out<=0;
   36475: out<=0;
   36476: out<=1;
   36477: out<=0;
   36478: out<=1;
   36479: out<=0;
   36480: out<=1;
   36481: out<=0;
   36482: out<=0;
   36483: out<=1;
   36484: out<=1;
   36485: out<=1;
   36486: out<=1;
   36487: out<=1;
   36488: out<=1;
   36489: out<=1;
   36490: out<=0;
   36491: out<=0;
   36492: out<=1;
   36493: out<=0;
   36494: out<=1;
   36495: out<=0;
   36496: out<=1;
   36497: out<=0;
   36498: out<=0;
   36499: out<=1;
   36500: out<=1;
   36501: out<=1;
   36502: out<=1;
   36503: out<=1;
   36504: out<=1;
   36505: out<=1;
   36506: out<=0;
   36507: out<=0;
   36508: out<=1;
   36509: out<=0;
   36510: out<=1;
   36511: out<=0;
   36512: out<=1;
   36513: out<=0;
   36514: out<=0;
   36515: out<=1;
   36516: out<=1;
   36517: out<=1;
   36518: out<=1;
   36519: out<=1;
   36520: out<=1;
   36521: out<=1;
   36522: out<=0;
   36523: out<=0;
   36524: out<=1;
   36525: out<=0;
   36526: out<=1;
   36527: out<=0;
   36528: out<=1;
   36529: out<=0;
   36530: out<=0;
   36531: out<=1;
   36532: out<=1;
   36533: out<=1;
   36534: out<=1;
   36535: out<=1;
   36536: out<=1;
   36537: out<=1;
   36538: out<=0;
   36539: out<=0;
   36540: out<=1;
   36541: out<=0;
   36542: out<=1;
   36543: out<=0;
   36544: out<=0;
   36545: out<=1;
   36546: out<=1;
   36547: out<=0;
   36548: out<=0;
   36549: out<=0;
   36550: out<=0;
   36551: out<=0;
   36552: out<=0;
   36553: out<=0;
   36554: out<=1;
   36555: out<=1;
   36556: out<=0;
   36557: out<=1;
   36558: out<=0;
   36559: out<=1;
   36560: out<=1;
   36561: out<=0;
   36562: out<=0;
   36563: out<=1;
   36564: out<=1;
   36565: out<=1;
   36566: out<=1;
   36567: out<=1;
   36568: out<=1;
   36569: out<=1;
   36570: out<=0;
   36571: out<=0;
   36572: out<=1;
   36573: out<=0;
   36574: out<=1;
   36575: out<=0;
   36576: out<=1;
   36577: out<=0;
   36578: out<=0;
   36579: out<=1;
   36580: out<=1;
   36581: out<=1;
   36582: out<=1;
   36583: out<=1;
   36584: out<=1;
   36585: out<=1;
   36586: out<=0;
   36587: out<=0;
   36588: out<=1;
   36589: out<=0;
   36590: out<=1;
   36591: out<=0;
   36592: out<=0;
   36593: out<=1;
   36594: out<=1;
   36595: out<=0;
   36596: out<=0;
   36597: out<=0;
   36598: out<=0;
   36599: out<=0;
   36600: out<=0;
   36601: out<=0;
   36602: out<=1;
   36603: out<=1;
   36604: out<=0;
   36605: out<=1;
   36606: out<=0;
   36607: out<=1;
   36608: out<=1;
   36609: out<=1;
   36610: out<=1;
   36611: out<=1;
   36612: out<=0;
   36613: out<=1;
   36614: out<=1;
   36615: out<=0;
   36616: out<=0;
   36617: out<=1;
   36618: out<=0;
   36619: out<=1;
   36620: out<=1;
   36621: out<=1;
   36622: out<=0;
   36623: out<=0;
   36624: out<=1;
   36625: out<=1;
   36626: out<=1;
   36627: out<=1;
   36628: out<=0;
   36629: out<=1;
   36630: out<=1;
   36631: out<=0;
   36632: out<=0;
   36633: out<=1;
   36634: out<=0;
   36635: out<=1;
   36636: out<=1;
   36637: out<=1;
   36638: out<=0;
   36639: out<=0;
   36640: out<=0;
   36641: out<=0;
   36642: out<=0;
   36643: out<=0;
   36644: out<=1;
   36645: out<=0;
   36646: out<=0;
   36647: out<=1;
   36648: out<=1;
   36649: out<=0;
   36650: out<=1;
   36651: out<=0;
   36652: out<=0;
   36653: out<=0;
   36654: out<=1;
   36655: out<=1;
   36656: out<=0;
   36657: out<=0;
   36658: out<=0;
   36659: out<=0;
   36660: out<=1;
   36661: out<=0;
   36662: out<=0;
   36663: out<=1;
   36664: out<=1;
   36665: out<=0;
   36666: out<=1;
   36667: out<=0;
   36668: out<=0;
   36669: out<=0;
   36670: out<=1;
   36671: out<=1;
   36672: out<=0;
   36673: out<=0;
   36674: out<=0;
   36675: out<=0;
   36676: out<=1;
   36677: out<=0;
   36678: out<=0;
   36679: out<=1;
   36680: out<=1;
   36681: out<=0;
   36682: out<=1;
   36683: out<=0;
   36684: out<=0;
   36685: out<=0;
   36686: out<=1;
   36687: out<=1;
   36688: out<=1;
   36689: out<=1;
   36690: out<=1;
   36691: out<=1;
   36692: out<=0;
   36693: out<=1;
   36694: out<=1;
   36695: out<=0;
   36696: out<=0;
   36697: out<=1;
   36698: out<=0;
   36699: out<=1;
   36700: out<=1;
   36701: out<=1;
   36702: out<=0;
   36703: out<=0;
   36704: out<=0;
   36705: out<=0;
   36706: out<=0;
   36707: out<=0;
   36708: out<=1;
   36709: out<=0;
   36710: out<=0;
   36711: out<=1;
   36712: out<=1;
   36713: out<=0;
   36714: out<=1;
   36715: out<=0;
   36716: out<=0;
   36717: out<=0;
   36718: out<=1;
   36719: out<=1;
   36720: out<=1;
   36721: out<=1;
   36722: out<=1;
   36723: out<=1;
   36724: out<=0;
   36725: out<=1;
   36726: out<=1;
   36727: out<=0;
   36728: out<=0;
   36729: out<=1;
   36730: out<=0;
   36731: out<=1;
   36732: out<=1;
   36733: out<=1;
   36734: out<=0;
   36735: out<=0;
   36736: out<=1;
   36737: out<=1;
   36738: out<=1;
   36739: out<=1;
   36740: out<=0;
   36741: out<=1;
   36742: out<=1;
   36743: out<=0;
   36744: out<=0;
   36745: out<=1;
   36746: out<=0;
   36747: out<=1;
   36748: out<=1;
   36749: out<=1;
   36750: out<=0;
   36751: out<=0;
   36752: out<=0;
   36753: out<=0;
   36754: out<=0;
   36755: out<=0;
   36756: out<=1;
   36757: out<=0;
   36758: out<=0;
   36759: out<=1;
   36760: out<=1;
   36761: out<=0;
   36762: out<=1;
   36763: out<=0;
   36764: out<=0;
   36765: out<=0;
   36766: out<=1;
   36767: out<=1;
   36768: out<=0;
   36769: out<=0;
   36770: out<=0;
   36771: out<=0;
   36772: out<=1;
   36773: out<=0;
   36774: out<=0;
   36775: out<=1;
   36776: out<=1;
   36777: out<=0;
   36778: out<=1;
   36779: out<=0;
   36780: out<=0;
   36781: out<=0;
   36782: out<=1;
   36783: out<=1;
   36784: out<=1;
   36785: out<=1;
   36786: out<=1;
   36787: out<=1;
   36788: out<=0;
   36789: out<=1;
   36790: out<=1;
   36791: out<=0;
   36792: out<=0;
   36793: out<=1;
   36794: out<=0;
   36795: out<=1;
   36796: out<=1;
   36797: out<=1;
   36798: out<=0;
   36799: out<=0;
   36800: out<=0;
   36801: out<=0;
   36802: out<=0;
   36803: out<=0;
   36804: out<=1;
   36805: out<=0;
   36806: out<=0;
   36807: out<=1;
   36808: out<=1;
   36809: out<=0;
   36810: out<=1;
   36811: out<=0;
   36812: out<=0;
   36813: out<=0;
   36814: out<=1;
   36815: out<=1;
   36816: out<=0;
   36817: out<=0;
   36818: out<=0;
   36819: out<=0;
   36820: out<=1;
   36821: out<=0;
   36822: out<=0;
   36823: out<=1;
   36824: out<=1;
   36825: out<=0;
   36826: out<=1;
   36827: out<=0;
   36828: out<=0;
   36829: out<=0;
   36830: out<=1;
   36831: out<=1;
   36832: out<=0;
   36833: out<=0;
   36834: out<=0;
   36835: out<=0;
   36836: out<=1;
   36837: out<=0;
   36838: out<=0;
   36839: out<=1;
   36840: out<=1;
   36841: out<=0;
   36842: out<=1;
   36843: out<=0;
   36844: out<=0;
   36845: out<=0;
   36846: out<=1;
   36847: out<=1;
   36848: out<=0;
   36849: out<=0;
   36850: out<=0;
   36851: out<=0;
   36852: out<=1;
   36853: out<=0;
   36854: out<=0;
   36855: out<=1;
   36856: out<=1;
   36857: out<=0;
   36858: out<=1;
   36859: out<=0;
   36860: out<=0;
   36861: out<=0;
   36862: out<=1;
   36863: out<=1;
   36864: out<=1;
   36865: out<=0;
   36866: out<=0;
   36867: out<=1;
   36868: out<=0;
   36869: out<=0;
   36870: out<=0;
   36871: out<=0;
   36872: out<=1;
   36873: out<=1;
   36874: out<=0;
   36875: out<=0;
   36876: out<=0;
   36877: out<=1;
   36878: out<=0;
   36879: out<=1;
   36880: out<=0;
   36881: out<=1;
   36882: out<=1;
   36883: out<=0;
   36884: out<=1;
   36885: out<=1;
   36886: out<=1;
   36887: out<=1;
   36888: out<=0;
   36889: out<=0;
   36890: out<=1;
   36891: out<=1;
   36892: out<=1;
   36893: out<=0;
   36894: out<=1;
   36895: out<=0;
   36896: out<=0;
   36897: out<=1;
   36898: out<=1;
   36899: out<=0;
   36900: out<=1;
   36901: out<=1;
   36902: out<=1;
   36903: out<=1;
   36904: out<=0;
   36905: out<=0;
   36906: out<=1;
   36907: out<=1;
   36908: out<=1;
   36909: out<=0;
   36910: out<=1;
   36911: out<=0;
   36912: out<=1;
   36913: out<=0;
   36914: out<=0;
   36915: out<=1;
   36916: out<=0;
   36917: out<=0;
   36918: out<=0;
   36919: out<=0;
   36920: out<=1;
   36921: out<=1;
   36922: out<=0;
   36923: out<=0;
   36924: out<=0;
   36925: out<=1;
   36926: out<=0;
   36927: out<=1;
   36928: out<=1;
   36929: out<=0;
   36930: out<=0;
   36931: out<=1;
   36932: out<=0;
   36933: out<=0;
   36934: out<=0;
   36935: out<=0;
   36936: out<=1;
   36937: out<=1;
   36938: out<=0;
   36939: out<=0;
   36940: out<=0;
   36941: out<=1;
   36942: out<=0;
   36943: out<=1;
   36944: out<=1;
   36945: out<=0;
   36946: out<=0;
   36947: out<=1;
   36948: out<=0;
   36949: out<=0;
   36950: out<=0;
   36951: out<=0;
   36952: out<=1;
   36953: out<=1;
   36954: out<=0;
   36955: out<=0;
   36956: out<=0;
   36957: out<=1;
   36958: out<=0;
   36959: out<=1;
   36960: out<=1;
   36961: out<=0;
   36962: out<=0;
   36963: out<=1;
   36964: out<=0;
   36965: out<=0;
   36966: out<=0;
   36967: out<=0;
   36968: out<=1;
   36969: out<=1;
   36970: out<=0;
   36971: out<=0;
   36972: out<=0;
   36973: out<=1;
   36974: out<=0;
   36975: out<=1;
   36976: out<=1;
   36977: out<=0;
   36978: out<=0;
   36979: out<=1;
   36980: out<=0;
   36981: out<=0;
   36982: out<=0;
   36983: out<=0;
   36984: out<=1;
   36985: out<=1;
   36986: out<=0;
   36987: out<=0;
   36988: out<=0;
   36989: out<=1;
   36990: out<=0;
   36991: out<=1;
   36992: out<=0;
   36993: out<=1;
   36994: out<=1;
   36995: out<=0;
   36996: out<=1;
   36997: out<=1;
   36998: out<=1;
   36999: out<=1;
   37000: out<=0;
   37001: out<=0;
   37002: out<=1;
   37003: out<=1;
   37004: out<=1;
   37005: out<=0;
   37006: out<=1;
   37007: out<=0;
   37008: out<=0;
   37009: out<=1;
   37010: out<=1;
   37011: out<=0;
   37012: out<=1;
   37013: out<=1;
   37014: out<=1;
   37015: out<=1;
   37016: out<=0;
   37017: out<=0;
   37018: out<=1;
   37019: out<=1;
   37020: out<=1;
   37021: out<=0;
   37022: out<=1;
   37023: out<=0;
   37024: out<=1;
   37025: out<=0;
   37026: out<=0;
   37027: out<=1;
   37028: out<=0;
   37029: out<=0;
   37030: out<=0;
   37031: out<=0;
   37032: out<=1;
   37033: out<=1;
   37034: out<=0;
   37035: out<=0;
   37036: out<=0;
   37037: out<=1;
   37038: out<=0;
   37039: out<=1;
   37040: out<=1;
   37041: out<=0;
   37042: out<=0;
   37043: out<=1;
   37044: out<=0;
   37045: out<=0;
   37046: out<=0;
   37047: out<=0;
   37048: out<=1;
   37049: out<=1;
   37050: out<=0;
   37051: out<=0;
   37052: out<=0;
   37053: out<=1;
   37054: out<=0;
   37055: out<=1;
   37056: out<=0;
   37057: out<=1;
   37058: out<=1;
   37059: out<=0;
   37060: out<=1;
   37061: out<=1;
   37062: out<=1;
   37063: out<=1;
   37064: out<=0;
   37065: out<=0;
   37066: out<=1;
   37067: out<=1;
   37068: out<=1;
   37069: out<=0;
   37070: out<=1;
   37071: out<=0;
   37072: out<=1;
   37073: out<=0;
   37074: out<=0;
   37075: out<=1;
   37076: out<=0;
   37077: out<=0;
   37078: out<=0;
   37079: out<=0;
   37080: out<=1;
   37081: out<=1;
   37082: out<=0;
   37083: out<=0;
   37084: out<=0;
   37085: out<=1;
   37086: out<=0;
   37087: out<=1;
   37088: out<=0;
   37089: out<=1;
   37090: out<=1;
   37091: out<=0;
   37092: out<=1;
   37093: out<=1;
   37094: out<=1;
   37095: out<=1;
   37096: out<=0;
   37097: out<=0;
   37098: out<=1;
   37099: out<=1;
   37100: out<=1;
   37101: out<=0;
   37102: out<=1;
   37103: out<=0;
   37104: out<=1;
   37105: out<=0;
   37106: out<=0;
   37107: out<=1;
   37108: out<=0;
   37109: out<=0;
   37110: out<=0;
   37111: out<=0;
   37112: out<=1;
   37113: out<=1;
   37114: out<=0;
   37115: out<=0;
   37116: out<=0;
   37117: out<=1;
   37118: out<=0;
   37119: out<=1;
   37120: out<=1;
   37121: out<=1;
   37122: out<=1;
   37123: out<=1;
   37124: out<=1;
   37125: out<=0;
   37126: out<=0;
   37127: out<=1;
   37128: out<=0;
   37129: out<=1;
   37130: out<=0;
   37131: out<=1;
   37132: out<=0;
   37133: out<=0;
   37134: out<=1;
   37135: out<=1;
   37136: out<=1;
   37137: out<=1;
   37138: out<=1;
   37139: out<=1;
   37140: out<=1;
   37141: out<=0;
   37142: out<=0;
   37143: out<=1;
   37144: out<=0;
   37145: out<=1;
   37146: out<=0;
   37147: out<=1;
   37148: out<=0;
   37149: out<=0;
   37150: out<=1;
   37151: out<=1;
   37152: out<=1;
   37153: out<=1;
   37154: out<=1;
   37155: out<=1;
   37156: out<=1;
   37157: out<=0;
   37158: out<=0;
   37159: out<=1;
   37160: out<=0;
   37161: out<=1;
   37162: out<=0;
   37163: out<=1;
   37164: out<=0;
   37165: out<=0;
   37166: out<=1;
   37167: out<=1;
   37168: out<=1;
   37169: out<=1;
   37170: out<=1;
   37171: out<=1;
   37172: out<=1;
   37173: out<=0;
   37174: out<=0;
   37175: out<=1;
   37176: out<=0;
   37177: out<=1;
   37178: out<=0;
   37179: out<=1;
   37180: out<=0;
   37181: out<=0;
   37182: out<=1;
   37183: out<=1;
   37184: out<=1;
   37185: out<=1;
   37186: out<=1;
   37187: out<=1;
   37188: out<=1;
   37189: out<=0;
   37190: out<=0;
   37191: out<=1;
   37192: out<=0;
   37193: out<=1;
   37194: out<=0;
   37195: out<=1;
   37196: out<=0;
   37197: out<=0;
   37198: out<=1;
   37199: out<=1;
   37200: out<=0;
   37201: out<=0;
   37202: out<=0;
   37203: out<=0;
   37204: out<=0;
   37205: out<=1;
   37206: out<=1;
   37207: out<=0;
   37208: out<=1;
   37209: out<=0;
   37210: out<=1;
   37211: out<=0;
   37212: out<=1;
   37213: out<=1;
   37214: out<=0;
   37215: out<=0;
   37216: out<=0;
   37217: out<=0;
   37218: out<=0;
   37219: out<=0;
   37220: out<=0;
   37221: out<=1;
   37222: out<=1;
   37223: out<=0;
   37224: out<=1;
   37225: out<=0;
   37226: out<=1;
   37227: out<=0;
   37228: out<=1;
   37229: out<=1;
   37230: out<=0;
   37231: out<=0;
   37232: out<=1;
   37233: out<=1;
   37234: out<=1;
   37235: out<=1;
   37236: out<=1;
   37237: out<=0;
   37238: out<=0;
   37239: out<=1;
   37240: out<=0;
   37241: out<=1;
   37242: out<=0;
   37243: out<=1;
   37244: out<=0;
   37245: out<=0;
   37246: out<=1;
   37247: out<=1;
   37248: out<=0;
   37249: out<=0;
   37250: out<=0;
   37251: out<=0;
   37252: out<=0;
   37253: out<=1;
   37254: out<=1;
   37255: out<=0;
   37256: out<=1;
   37257: out<=0;
   37258: out<=1;
   37259: out<=0;
   37260: out<=1;
   37261: out<=1;
   37262: out<=0;
   37263: out<=0;
   37264: out<=1;
   37265: out<=1;
   37266: out<=1;
   37267: out<=1;
   37268: out<=1;
   37269: out<=0;
   37270: out<=0;
   37271: out<=1;
   37272: out<=0;
   37273: out<=1;
   37274: out<=0;
   37275: out<=1;
   37276: out<=0;
   37277: out<=0;
   37278: out<=1;
   37279: out<=1;
   37280: out<=0;
   37281: out<=0;
   37282: out<=0;
   37283: out<=0;
   37284: out<=0;
   37285: out<=1;
   37286: out<=1;
   37287: out<=0;
   37288: out<=1;
   37289: out<=0;
   37290: out<=1;
   37291: out<=0;
   37292: out<=1;
   37293: out<=1;
   37294: out<=0;
   37295: out<=0;
   37296: out<=1;
   37297: out<=1;
   37298: out<=1;
   37299: out<=1;
   37300: out<=1;
   37301: out<=0;
   37302: out<=0;
   37303: out<=1;
   37304: out<=0;
   37305: out<=1;
   37306: out<=0;
   37307: out<=1;
   37308: out<=0;
   37309: out<=0;
   37310: out<=1;
   37311: out<=1;
   37312: out<=0;
   37313: out<=0;
   37314: out<=0;
   37315: out<=0;
   37316: out<=0;
   37317: out<=1;
   37318: out<=1;
   37319: out<=0;
   37320: out<=1;
   37321: out<=0;
   37322: out<=1;
   37323: out<=0;
   37324: out<=1;
   37325: out<=1;
   37326: out<=0;
   37327: out<=0;
   37328: out<=0;
   37329: out<=0;
   37330: out<=0;
   37331: out<=0;
   37332: out<=0;
   37333: out<=1;
   37334: out<=1;
   37335: out<=0;
   37336: out<=1;
   37337: out<=0;
   37338: out<=1;
   37339: out<=0;
   37340: out<=1;
   37341: out<=1;
   37342: out<=0;
   37343: out<=0;
   37344: out<=1;
   37345: out<=1;
   37346: out<=1;
   37347: out<=1;
   37348: out<=1;
   37349: out<=0;
   37350: out<=0;
   37351: out<=1;
   37352: out<=0;
   37353: out<=1;
   37354: out<=0;
   37355: out<=1;
   37356: out<=0;
   37357: out<=0;
   37358: out<=1;
   37359: out<=1;
   37360: out<=1;
   37361: out<=1;
   37362: out<=1;
   37363: out<=1;
   37364: out<=1;
   37365: out<=0;
   37366: out<=0;
   37367: out<=1;
   37368: out<=0;
   37369: out<=1;
   37370: out<=0;
   37371: out<=1;
   37372: out<=0;
   37373: out<=0;
   37374: out<=1;
   37375: out<=1;
   37376: out<=1;
   37377: out<=1;
   37378: out<=0;
   37379: out<=0;
   37380: out<=1;
   37381: out<=0;
   37382: out<=1;
   37383: out<=0;
   37384: out<=1;
   37385: out<=0;
   37386: out<=0;
   37387: out<=1;
   37388: out<=1;
   37389: out<=1;
   37390: out<=1;
   37391: out<=1;
   37392: out<=1;
   37393: out<=1;
   37394: out<=0;
   37395: out<=0;
   37396: out<=1;
   37397: out<=0;
   37398: out<=1;
   37399: out<=0;
   37400: out<=1;
   37401: out<=0;
   37402: out<=0;
   37403: out<=1;
   37404: out<=1;
   37405: out<=1;
   37406: out<=1;
   37407: out<=1;
   37408: out<=0;
   37409: out<=0;
   37410: out<=1;
   37411: out<=1;
   37412: out<=0;
   37413: out<=1;
   37414: out<=0;
   37415: out<=1;
   37416: out<=0;
   37417: out<=1;
   37418: out<=1;
   37419: out<=0;
   37420: out<=0;
   37421: out<=0;
   37422: out<=0;
   37423: out<=0;
   37424: out<=0;
   37425: out<=0;
   37426: out<=1;
   37427: out<=1;
   37428: out<=0;
   37429: out<=1;
   37430: out<=0;
   37431: out<=1;
   37432: out<=0;
   37433: out<=1;
   37434: out<=1;
   37435: out<=0;
   37436: out<=0;
   37437: out<=0;
   37438: out<=0;
   37439: out<=0;
   37440: out<=1;
   37441: out<=1;
   37442: out<=0;
   37443: out<=0;
   37444: out<=1;
   37445: out<=0;
   37446: out<=1;
   37447: out<=0;
   37448: out<=1;
   37449: out<=0;
   37450: out<=0;
   37451: out<=1;
   37452: out<=1;
   37453: out<=1;
   37454: out<=1;
   37455: out<=1;
   37456: out<=0;
   37457: out<=0;
   37458: out<=1;
   37459: out<=1;
   37460: out<=0;
   37461: out<=1;
   37462: out<=0;
   37463: out<=1;
   37464: out<=0;
   37465: out<=1;
   37466: out<=1;
   37467: out<=0;
   37468: out<=0;
   37469: out<=0;
   37470: out<=0;
   37471: out<=0;
   37472: out<=1;
   37473: out<=1;
   37474: out<=0;
   37475: out<=0;
   37476: out<=1;
   37477: out<=0;
   37478: out<=1;
   37479: out<=0;
   37480: out<=1;
   37481: out<=0;
   37482: out<=0;
   37483: out<=1;
   37484: out<=1;
   37485: out<=1;
   37486: out<=1;
   37487: out<=1;
   37488: out<=0;
   37489: out<=0;
   37490: out<=1;
   37491: out<=1;
   37492: out<=0;
   37493: out<=1;
   37494: out<=0;
   37495: out<=1;
   37496: out<=0;
   37497: out<=1;
   37498: out<=1;
   37499: out<=0;
   37500: out<=0;
   37501: out<=0;
   37502: out<=0;
   37503: out<=0;
   37504: out<=0;
   37505: out<=0;
   37506: out<=1;
   37507: out<=1;
   37508: out<=0;
   37509: out<=1;
   37510: out<=0;
   37511: out<=1;
   37512: out<=0;
   37513: out<=1;
   37514: out<=1;
   37515: out<=0;
   37516: out<=0;
   37517: out<=0;
   37518: out<=0;
   37519: out<=0;
   37520: out<=1;
   37521: out<=1;
   37522: out<=0;
   37523: out<=0;
   37524: out<=1;
   37525: out<=0;
   37526: out<=1;
   37527: out<=0;
   37528: out<=1;
   37529: out<=0;
   37530: out<=0;
   37531: out<=1;
   37532: out<=1;
   37533: out<=1;
   37534: out<=1;
   37535: out<=1;
   37536: out<=1;
   37537: out<=1;
   37538: out<=0;
   37539: out<=0;
   37540: out<=1;
   37541: out<=0;
   37542: out<=1;
   37543: out<=0;
   37544: out<=1;
   37545: out<=0;
   37546: out<=0;
   37547: out<=1;
   37548: out<=1;
   37549: out<=1;
   37550: out<=1;
   37551: out<=1;
   37552: out<=0;
   37553: out<=0;
   37554: out<=1;
   37555: out<=1;
   37556: out<=0;
   37557: out<=1;
   37558: out<=0;
   37559: out<=1;
   37560: out<=0;
   37561: out<=1;
   37562: out<=1;
   37563: out<=0;
   37564: out<=0;
   37565: out<=0;
   37566: out<=0;
   37567: out<=0;
   37568: out<=0;
   37569: out<=0;
   37570: out<=1;
   37571: out<=1;
   37572: out<=0;
   37573: out<=1;
   37574: out<=0;
   37575: out<=1;
   37576: out<=0;
   37577: out<=1;
   37578: out<=1;
   37579: out<=0;
   37580: out<=0;
   37581: out<=0;
   37582: out<=0;
   37583: out<=0;
   37584: out<=0;
   37585: out<=0;
   37586: out<=1;
   37587: out<=1;
   37588: out<=0;
   37589: out<=1;
   37590: out<=0;
   37591: out<=1;
   37592: out<=0;
   37593: out<=1;
   37594: out<=1;
   37595: out<=0;
   37596: out<=0;
   37597: out<=0;
   37598: out<=0;
   37599: out<=0;
   37600: out<=0;
   37601: out<=0;
   37602: out<=1;
   37603: out<=1;
   37604: out<=0;
   37605: out<=1;
   37606: out<=0;
   37607: out<=1;
   37608: out<=0;
   37609: out<=1;
   37610: out<=1;
   37611: out<=0;
   37612: out<=0;
   37613: out<=0;
   37614: out<=0;
   37615: out<=0;
   37616: out<=0;
   37617: out<=0;
   37618: out<=1;
   37619: out<=1;
   37620: out<=0;
   37621: out<=1;
   37622: out<=0;
   37623: out<=1;
   37624: out<=0;
   37625: out<=1;
   37626: out<=1;
   37627: out<=0;
   37628: out<=0;
   37629: out<=0;
   37630: out<=0;
   37631: out<=0;
   37632: out<=1;
   37633: out<=0;
   37634: out<=1;
   37635: out<=0;
   37636: out<=0;
   37637: out<=0;
   37638: out<=1;
   37639: out<=1;
   37640: out<=0;
   37641: out<=0;
   37642: out<=0;
   37643: out<=0;
   37644: out<=1;
   37645: out<=0;
   37646: out<=0;
   37647: out<=1;
   37648: out<=0;
   37649: out<=1;
   37650: out<=0;
   37651: out<=1;
   37652: out<=1;
   37653: out<=1;
   37654: out<=0;
   37655: out<=0;
   37656: out<=1;
   37657: out<=1;
   37658: out<=1;
   37659: out<=1;
   37660: out<=0;
   37661: out<=1;
   37662: out<=1;
   37663: out<=0;
   37664: out<=1;
   37665: out<=0;
   37666: out<=1;
   37667: out<=0;
   37668: out<=0;
   37669: out<=0;
   37670: out<=1;
   37671: out<=1;
   37672: out<=0;
   37673: out<=0;
   37674: out<=0;
   37675: out<=0;
   37676: out<=1;
   37677: out<=0;
   37678: out<=0;
   37679: out<=1;
   37680: out<=0;
   37681: out<=1;
   37682: out<=0;
   37683: out<=1;
   37684: out<=1;
   37685: out<=1;
   37686: out<=0;
   37687: out<=0;
   37688: out<=1;
   37689: out<=1;
   37690: out<=1;
   37691: out<=1;
   37692: out<=0;
   37693: out<=1;
   37694: out<=1;
   37695: out<=0;
   37696: out<=1;
   37697: out<=0;
   37698: out<=1;
   37699: out<=0;
   37700: out<=0;
   37701: out<=0;
   37702: out<=1;
   37703: out<=1;
   37704: out<=0;
   37705: out<=0;
   37706: out<=0;
   37707: out<=0;
   37708: out<=1;
   37709: out<=0;
   37710: out<=0;
   37711: out<=1;
   37712: out<=1;
   37713: out<=0;
   37714: out<=1;
   37715: out<=0;
   37716: out<=0;
   37717: out<=0;
   37718: out<=1;
   37719: out<=1;
   37720: out<=0;
   37721: out<=0;
   37722: out<=0;
   37723: out<=0;
   37724: out<=1;
   37725: out<=0;
   37726: out<=0;
   37727: out<=1;
   37728: out<=0;
   37729: out<=1;
   37730: out<=0;
   37731: out<=1;
   37732: out<=1;
   37733: out<=1;
   37734: out<=0;
   37735: out<=0;
   37736: out<=1;
   37737: out<=1;
   37738: out<=1;
   37739: out<=1;
   37740: out<=0;
   37741: out<=1;
   37742: out<=1;
   37743: out<=0;
   37744: out<=0;
   37745: out<=1;
   37746: out<=0;
   37747: out<=1;
   37748: out<=1;
   37749: out<=1;
   37750: out<=0;
   37751: out<=0;
   37752: out<=1;
   37753: out<=1;
   37754: out<=1;
   37755: out<=1;
   37756: out<=0;
   37757: out<=1;
   37758: out<=1;
   37759: out<=0;
   37760: out<=0;
   37761: out<=1;
   37762: out<=0;
   37763: out<=1;
   37764: out<=1;
   37765: out<=1;
   37766: out<=0;
   37767: out<=0;
   37768: out<=1;
   37769: out<=1;
   37770: out<=1;
   37771: out<=1;
   37772: out<=0;
   37773: out<=1;
   37774: out<=1;
   37775: out<=0;
   37776: out<=0;
   37777: out<=1;
   37778: out<=0;
   37779: out<=1;
   37780: out<=1;
   37781: out<=1;
   37782: out<=0;
   37783: out<=0;
   37784: out<=1;
   37785: out<=1;
   37786: out<=1;
   37787: out<=1;
   37788: out<=0;
   37789: out<=1;
   37790: out<=1;
   37791: out<=0;
   37792: out<=0;
   37793: out<=1;
   37794: out<=0;
   37795: out<=1;
   37796: out<=1;
   37797: out<=1;
   37798: out<=0;
   37799: out<=0;
   37800: out<=1;
   37801: out<=1;
   37802: out<=1;
   37803: out<=1;
   37804: out<=0;
   37805: out<=1;
   37806: out<=1;
   37807: out<=0;
   37808: out<=0;
   37809: out<=1;
   37810: out<=0;
   37811: out<=1;
   37812: out<=1;
   37813: out<=1;
   37814: out<=0;
   37815: out<=0;
   37816: out<=1;
   37817: out<=1;
   37818: out<=1;
   37819: out<=1;
   37820: out<=0;
   37821: out<=1;
   37822: out<=1;
   37823: out<=0;
   37824: out<=0;
   37825: out<=1;
   37826: out<=0;
   37827: out<=1;
   37828: out<=1;
   37829: out<=1;
   37830: out<=0;
   37831: out<=0;
   37832: out<=1;
   37833: out<=1;
   37834: out<=1;
   37835: out<=1;
   37836: out<=0;
   37837: out<=1;
   37838: out<=1;
   37839: out<=0;
   37840: out<=1;
   37841: out<=0;
   37842: out<=1;
   37843: out<=0;
   37844: out<=0;
   37845: out<=0;
   37846: out<=1;
   37847: out<=1;
   37848: out<=0;
   37849: out<=0;
   37850: out<=0;
   37851: out<=0;
   37852: out<=1;
   37853: out<=0;
   37854: out<=0;
   37855: out<=1;
   37856: out<=1;
   37857: out<=0;
   37858: out<=1;
   37859: out<=0;
   37860: out<=0;
   37861: out<=0;
   37862: out<=1;
   37863: out<=1;
   37864: out<=0;
   37865: out<=0;
   37866: out<=0;
   37867: out<=0;
   37868: out<=1;
   37869: out<=0;
   37870: out<=0;
   37871: out<=1;
   37872: out<=0;
   37873: out<=1;
   37874: out<=0;
   37875: out<=1;
   37876: out<=1;
   37877: out<=1;
   37878: out<=0;
   37879: out<=0;
   37880: out<=1;
   37881: out<=1;
   37882: out<=1;
   37883: out<=1;
   37884: out<=0;
   37885: out<=1;
   37886: out<=1;
   37887: out<=0;
   37888: out<=1;
   37889: out<=1;
   37890: out<=1;
   37891: out<=1;
   37892: out<=0;
   37893: out<=1;
   37894: out<=1;
   37895: out<=0;
   37896: out<=1;
   37897: out<=0;
   37898: out<=1;
   37899: out<=0;
   37900: out<=0;
   37901: out<=0;
   37902: out<=1;
   37903: out<=1;
   37904: out<=0;
   37905: out<=0;
   37906: out<=0;
   37907: out<=0;
   37908: out<=1;
   37909: out<=0;
   37910: out<=0;
   37911: out<=1;
   37912: out<=0;
   37913: out<=1;
   37914: out<=0;
   37915: out<=1;
   37916: out<=1;
   37917: out<=1;
   37918: out<=0;
   37919: out<=0;
   37920: out<=0;
   37921: out<=0;
   37922: out<=0;
   37923: out<=0;
   37924: out<=1;
   37925: out<=0;
   37926: out<=0;
   37927: out<=1;
   37928: out<=0;
   37929: out<=1;
   37930: out<=0;
   37931: out<=1;
   37932: out<=1;
   37933: out<=1;
   37934: out<=0;
   37935: out<=0;
   37936: out<=1;
   37937: out<=1;
   37938: out<=1;
   37939: out<=1;
   37940: out<=0;
   37941: out<=1;
   37942: out<=1;
   37943: out<=0;
   37944: out<=1;
   37945: out<=0;
   37946: out<=1;
   37947: out<=0;
   37948: out<=0;
   37949: out<=0;
   37950: out<=1;
   37951: out<=1;
   37952: out<=1;
   37953: out<=1;
   37954: out<=1;
   37955: out<=1;
   37956: out<=0;
   37957: out<=1;
   37958: out<=1;
   37959: out<=0;
   37960: out<=1;
   37961: out<=0;
   37962: out<=1;
   37963: out<=0;
   37964: out<=0;
   37965: out<=0;
   37966: out<=1;
   37967: out<=1;
   37968: out<=1;
   37969: out<=1;
   37970: out<=1;
   37971: out<=1;
   37972: out<=0;
   37973: out<=1;
   37974: out<=1;
   37975: out<=0;
   37976: out<=1;
   37977: out<=0;
   37978: out<=1;
   37979: out<=0;
   37980: out<=0;
   37981: out<=0;
   37982: out<=1;
   37983: out<=1;
   37984: out<=1;
   37985: out<=1;
   37986: out<=1;
   37987: out<=1;
   37988: out<=0;
   37989: out<=1;
   37990: out<=1;
   37991: out<=0;
   37992: out<=1;
   37993: out<=0;
   37994: out<=1;
   37995: out<=0;
   37996: out<=0;
   37997: out<=0;
   37998: out<=1;
   37999: out<=1;
   38000: out<=1;
   38001: out<=1;
   38002: out<=1;
   38003: out<=1;
   38004: out<=0;
   38005: out<=1;
   38006: out<=1;
   38007: out<=0;
   38008: out<=1;
   38009: out<=0;
   38010: out<=1;
   38011: out<=0;
   38012: out<=0;
   38013: out<=0;
   38014: out<=1;
   38015: out<=1;
   38016: out<=0;
   38017: out<=0;
   38018: out<=0;
   38019: out<=0;
   38020: out<=1;
   38021: out<=0;
   38022: out<=0;
   38023: out<=1;
   38024: out<=0;
   38025: out<=1;
   38026: out<=0;
   38027: out<=1;
   38028: out<=1;
   38029: out<=1;
   38030: out<=0;
   38031: out<=0;
   38032: out<=0;
   38033: out<=0;
   38034: out<=0;
   38035: out<=0;
   38036: out<=1;
   38037: out<=0;
   38038: out<=0;
   38039: out<=1;
   38040: out<=0;
   38041: out<=1;
   38042: out<=0;
   38043: out<=1;
   38044: out<=1;
   38045: out<=1;
   38046: out<=0;
   38047: out<=0;
   38048: out<=1;
   38049: out<=1;
   38050: out<=1;
   38051: out<=1;
   38052: out<=0;
   38053: out<=1;
   38054: out<=1;
   38055: out<=0;
   38056: out<=1;
   38057: out<=0;
   38058: out<=1;
   38059: out<=0;
   38060: out<=0;
   38061: out<=0;
   38062: out<=1;
   38063: out<=1;
   38064: out<=1;
   38065: out<=1;
   38066: out<=1;
   38067: out<=1;
   38068: out<=0;
   38069: out<=1;
   38070: out<=1;
   38071: out<=0;
   38072: out<=1;
   38073: out<=0;
   38074: out<=1;
   38075: out<=0;
   38076: out<=0;
   38077: out<=0;
   38078: out<=1;
   38079: out<=1;
   38080: out<=0;
   38081: out<=0;
   38082: out<=0;
   38083: out<=0;
   38084: out<=1;
   38085: out<=0;
   38086: out<=0;
   38087: out<=1;
   38088: out<=0;
   38089: out<=1;
   38090: out<=0;
   38091: out<=1;
   38092: out<=1;
   38093: out<=1;
   38094: out<=0;
   38095: out<=0;
   38096: out<=1;
   38097: out<=1;
   38098: out<=1;
   38099: out<=1;
   38100: out<=0;
   38101: out<=1;
   38102: out<=1;
   38103: out<=0;
   38104: out<=1;
   38105: out<=0;
   38106: out<=1;
   38107: out<=0;
   38108: out<=0;
   38109: out<=0;
   38110: out<=1;
   38111: out<=1;
   38112: out<=0;
   38113: out<=0;
   38114: out<=0;
   38115: out<=0;
   38116: out<=1;
   38117: out<=0;
   38118: out<=0;
   38119: out<=1;
   38120: out<=0;
   38121: out<=1;
   38122: out<=0;
   38123: out<=1;
   38124: out<=1;
   38125: out<=1;
   38126: out<=0;
   38127: out<=0;
   38128: out<=1;
   38129: out<=1;
   38130: out<=1;
   38131: out<=1;
   38132: out<=0;
   38133: out<=1;
   38134: out<=1;
   38135: out<=0;
   38136: out<=1;
   38137: out<=0;
   38138: out<=1;
   38139: out<=0;
   38140: out<=0;
   38141: out<=0;
   38142: out<=1;
   38143: out<=1;
   38144: out<=0;
   38145: out<=1;
   38146: out<=1;
   38147: out<=0;
   38148: out<=0;
   38149: out<=0;
   38150: out<=0;
   38151: out<=0;
   38152: out<=1;
   38153: out<=1;
   38154: out<=0;
   38155: out<=0;
   38156: out<=1;
   38157: out<=0;
   38158: out<=1;
   38159: out<=0;
   38160: out<=0;
   38161: out<=1;
   38162: out<=1;
   38163: out<=0;
   38164: out<=0;
   38165: out<=0;
   38166: out<=0;
   38167: out<=0;
   38168: out<=1;
   38169: out<=1;
   38170: out<=0;
   38171: out<=0;
   38172: out<=1;
   38173: out<=0;
   38174: out<=1;
   38175: out<=0;
   38176: out<=0;
   38177: out<=1;
   38178: out<=1;
   38179: out<=0;
   38180: out<=0;
   38181: out<=0;
   38182: out<=0;
   38183: out<=0;
   38184: out<=1;
   38185: out<=1;
   38186: out<=0;
   38187: out<=0;
   38188: out<=1;
   38189: out<=0;
   38190: out<=1;
   38191: out<=0;
   38192: out<=0;
   38193: out<=1;
   38194: out<=1;
   38195: out<=0;
   38196: out<=0;
   38197: out<=0;
   38198: out<=0;
   38199: out<=0;
   38200: out<=1;
   38201: out<=1;
   38202: out<=0;
   38203: out<=0;
   38204: out<=1;
   38205: out<=0;
   38206: out<=1;
   38207: out<=0;
   38208: out<=0;
   38209: out<=1;
   38210: out<=1;
   38211: out<=0;
   38212: out<=0;
   38213: out<=0;
   38214: out<=0;
   38215: out<=0;
   38216: out<=1;
   38217: out<=1;
   38218: out<=0;
   38219: out<=0;
   38220: out<=1;
   38221: out<=0;
   38222: out<=1;
   38223: out<=0;
   38224: out<=1;
   38225: out<=0;
   38226: out<=0;
   38227: out<=1;
   38228: out<=1;
   38229: out<=1;
   38230: out<=1;
   38231: out<=1;
   38232: out<=0;
   38233: out<=0;
   38234: out<=1;
   38235: out<=1;
   38236: out<=0;
   38237: out<=1;
   38238: out<=0;
   38239: out<=1;
   38240: out<=1;
   38241: out<=0;
   38242: out<=0;
   38243: out<=1;
   38244: out<=1;
   38245: out<=1;
   38246: out<=1;
   38247: out<=1;
   38248: out<=0;
   38249: out<=0;
   38250: out<=1;
   38251: out<=1;
   38252: out<=0;
   38253: out<=1;
   38254: out<=0;
   38255: out<=1;
   38256: out<=0;
   38257: out<=1;
   38258: out<=1;
   38259: out<=0;
   38260: out<=0;
   38261: out<=0;
   38262: out<=0;
   38263: out<=0;
   38264: out<=1;
   38265: out<=1;
   38266: out<=0;
   38267: out<=0;
   38268: out<=1;
   38269: out<=0;
   38270: out<=1;
   38271: out<=0;
   38272: out<=1;
   38273: out<=0;
   38274: out<=0;
   38275: out<=1;
   38276: out<=1;
   38277: out<=1;
   38278: out<=1;
   38279: out<=1;
   38280: out<=0;
   38281: out<=0;
   38282: out<=1;
   38283: out<=1;
   38284: out<=0;
   38285: out<=1;
   38286: out<=0;
   38287: out<=1;
   38288: out<=0;
   38289: out<=1;
   38290: out<=1;
   38291: out<=0;
   38292: out<=0;
   38293: out<=0;
   38294: out<=0;
   38295: out<=0;
   38296: out<=1;
   38297: out<=1;
   38298: out<=0;
   38299: out<=0;
   38300: out<=1;
   38301: out<=0;
   38302: out<=1;
   38303: out<=0;
   38304: out<=1;
   38305: out<=0;
   38306: out<=0;
   38307: out<=1;
   38308: out<=1;
   38309: out<=1;
   38310: out<=1;
   38311: out<=1;
   38312: out<=0;
   38313: out<=0;
   38314: out<=1;
   38315: out<=1;
   38316: out<=0;
   38317: out<=1;
   38318: out<=0;
   38319: out<=1;
   38320: out<=0;
   38321: out<=1;
   38322: out<=1;
   38323: out<=0;
   38324: out<=0;
   38325: out<=0;
   38326: out<=0;
   38327: out<=0;
   38328: out<=1;
   38329: out<=1;
   38330: out<=0;
   38331: out<=0;
   38332: out<=1;
   38333: out<=0;
   38334: out<=1;
   38335: out<=0;
   38336: out<=1;
   38337: out<=0;
   38338: out<=0;
   38339: out<=1;
   38340: out<=1;
   38341: out<=1;
   38342: out<=1;
   38343: out<=1;
   38344: out<=0;
   38345: out<=0;
   38346: out<=1;
   38347: out<=1;
   38348: out<=0;
   38349: out<=1;
   38350: out<=0;
   38351: out<=1;
   38352: out<=1;
   38353: out<=0;
   38354: out<=0;
   38355: out<=1;
   38356: out<=1;
   38357: out<=1;
   38358: out<=1;
   38359: out<=1;
   38360: out<=0;
   38361: out<=0;
   38362: out<=1;
   38363: out<=1;
   38364: out<=0;
   38365: out<=1;
   38366: out<=0;
   38367: out<=1;
   38368: out<=0;
   38369: out<=1;
   38370: out<=1;
   38371: out<=0;
   38372: out<=0;
   38373: out<=0;
   38374: out<=0;
   38375: out<=0;
   38376: out<=1;
   38377: out<=1;
   38378: out<=0;
   38379: out<=0;
   38380: out<=1;
   38381: out<=0;
   38382: out<=1;
   38383: out<=0;
   38384: out<=0;
   38385: out<=1;
   38386: out<=1;
   38387: out<=0;
   38388: out<=0;
   38389: out<=0;
   38390: out<=0;
   38391: out<=0;
   38392: out<=1;
   38393: out<=1;
   38394: out<=0;
   38395: out<=0;
   38396: out<=1;
   38397: out<=0;
   38398: out<=1;
   38399: out<=0;
   38400: out<=0;
   38401: out<=1;
   38402: out<=0;
   38403: out<=1;
   38404: out<=0;
   38405: out<=0;
   38406: out<=1;
   38407: out<=1;
   38408: out<=0;
   38409: out<=0;
   38410: out<=0;
   38411: out<=0;
   38412: out<=0;
   38413: out<=1;
   38414: out<=1;
   38415: out<=0;
   38416: out<=0;
   38417: out<=1;
   38418: out<=0;
   38419: out<=1;
   38420: out<=0;
   38421: out<=0;
   38422: out<=1;
   38423: out<=1;
   38424: out<=0;
   38425: out<=0;
   38426: out<=0;
   38427: out<=0;
   38428: out<=0;
   38429: out<=1;
   38430: out<=1;
   38431: out<=0;
   38432: out<=1;
   38433: out<=0;
   38434: out<=1;
   38435: out<=0;
   38436: out<=1;
   38437: out<=1;
   38438: out<=0;
   38439: out<=0;
   38440: out<=1;
   38441: out<=1;
   38442: out<=1;
   38443: out<=1;
   38444: out<=1;
   38445: out<=0;
   38446: out<=0;
   38447: out<=1;
   38448: out<=1;
   38449: out<=0;
   38450: out<=1;
   38451: out<=0;
   38452: out<=1;
   38453: out<=1;
   38454: out<=0;
   38455: out<=0;
   38456: out<=1;
   38457: out<=1;
   38458: out<=1;
   38459: out<=1;
   38460: out<=1;
   38461: out<=0;
   38462: out<=0;
   38463: out<=1;
   38464: out<=0;
   38465: out<=1;
   38466: out<=0;
   38467: out<=1;
   38468: out<=0;
   38469: out<=0;
   38470: out<=1;
   38471: out<=1;
   38472: out<=0;
   38473: out<=0;
   38474: out<=0;
   38475: out<=0;
   38476: out<=0;
   38477: out<=1;
   38478: out<=1;
   38479: out<=0;
   38480: out<=1;
   38481: out<=0;
   38482: out<=1;
   38483: out<=0;
   38484: out<=1;
   38485: out<=1;
   38486: out<=0;
   38487: out<=0;
   38488: out<=1;
   38489: out<=1;
   38490: out<=1;
   38491: out<=1;
   38492: out<=1;
   38493: out<=0;
   38494: out<=0;
   38495: out<=1;
   38496: out<=0;
   38497: out<=1;
   38498: out<=0;
   38499: out<=1;
   38500: out<=0;
   38501: out<=0;
   38502: out<=1;
   38503: out<=1;
   38504: out<=0;
   38505: out<=0;
   38506: out<=0;
   38507: out<=0;
   38508: out<=0;
   38509: out<=1;
   38510: out<=1;
   38511: out<=0;
   38512: out<=1;
   38513: out<=0;
   38514: out<=1;
   38515: out<=0;
   38516: out<=1;
   38517: out<=1;
   38518: out<=0;
   38519: out<=0;
   38520: out<=1;
   38521: out<=1;
   38522: out<=1;
   38523: out<=1;
   38524: out<=1;
   38525: out<=0;
   38526: out<=0;
   38527: out<=1;
   38528: out<=1;
   38529: out<=0;
   38530: out<=1;
   38531: out<=0;
   38532: out<=1;
   38533: out<=1;
   38534: out<=0;
   38535: out<=0;
   38536: out<=1;
   38537: out<=1;
   38538: out<=1;
   38539: out<=1;
   38540: out<=1;
   38541: out<=0;
   38542: out<=0;
   38543: out<=1;
   38544: out<=0;
   38545: out<=1;
   38546: out<=0;
   38547: out<=1;
   38548: out<=0;
   38549: out<=0;
   38550: out<=1;
   38551: out<=1;
   38552: out<=0;
   38553: out<=0;
   38554: out<=0;
   38555: out<=0;
   38556: out<=0;
   38557: out<=1;
   38558: out<=1;
   38559: out<=0;
   38560: out<=0;
   38561: out<=1;
   38562: out<=0;
   38563: out<=1;
   38564: out<=0;
   38565: out<=0;
   38566: out<=1;
   38567: out<=1;
   38568: out<=0;
   38569: out<=0;
   38570: out<=0;
   38571: out<=0;
   38572: out<=0;
   38573: out<=1;
   38574: out<=1;
   38575: out<=0;
   38576: out<=1;
   38577: out<=0;
   38578: out<=1;
   38579: out<=0;
   38580: out<=1;
   38581: out<=1;
   38582: out<=0;
   38583: out<=0;
   38584: out<=1;
   38585: out<=1;
   38586: out<=1;
   38587: out<=1;
   38588: out<=1;
   38589: out<=0;
   38590: out<=0;
   38591: out<=1;
   38592: out<=1;
   38593: out<=0;
   38594: out<=1;
   38595: out<=0;
   38596: out<=1;
   38597: out<=1;
   38598: out<=0;
   38599: out<=0;
   38600: out<=1;
   38601: out<=1;
   38602: out<=1;
   38603: out<=1;
   38604: out<=1;
   38605: out<=0;
   38606: out<=0;
   38607: out<=1;
   38608: out<=1;
   38609: out<=0;
   38610: out<=1;
   38611: out<=0;
   38612: out<=1;
   38613: out<=1;
   38614: out<=0;
   38615: out<=0;
   38616: out<=1;
   38617: out<=1;
   38618: out<=1;
   38619: out<=1;
   38620: out<=1;
   38621: out<=0;
   38622: out<=0;
   38623: out<=1;
   38624: out<=1;
   38625: out<=0;
   38626: out<=1;
   38627: out<=0;
   38628: out<=1;
   38629: out<=1;
   38630: out<=0;
   38631: out<=0;
   38632: out<=1;
   38633: out<=1;
   38634: out<=1;
   38635: out<=1;
   38636: out<=1;
   38637: out<=0;
   38638: out<=0;
   38639: out<=1;
   38640: out<=1;
   38641: out<=0;
   38642: out<=1;
   38643: out<=0;
   38644: out<=1;
   38645: out<=1;
   38646: out<=0;
   38647: out<=0;
   38648: out<=1;
   38649: out<=1;
   38650: out<=1;
   38651: out<=1;
   38652: out<=1;
   38653: out<=0;
   38654: out<=0;
   38655: out<=1;
   38656: out<=1;
   38657: out<=1;
   38658: out<=0;
   38659: out<=0;
   38660: out<=0;
   38661: out<=1;
   38662: out<=0;
   38663: out<=1;
   38664: out<=0;
   38665: out<=1;
   38666: out<=1;
   38667: out<=0;
   38668: out<=1;
   38669: out<=1;
   38670: out<=1;
   38671: out<=1;
   38672: out<=0;
   38673: out<=0;
   38674: out<=1;
   38675: out<=1;
   38676: out<=1;
   38677: out<=0;
   38678: out<=1;
   38679: out<=0;
   38680: out<=1;
   38681: out<=0;
   38682: out<=0;
   38683: out<=1;
   38684: out<=0;
   38685: out<=0;
   38686: out<=0;
   38687: out<=0;
   38688: out<=1;
   38689: out<=1;
   38690: out<=0;
   38691: out<=0;
   38692: out<=0;
   38693: out<=1;
   38694: out<=0;
   38695: out<=1;
   38696: out<=0;
   38697: out<=1;
   38698: out<=1;
   38699: out<=0;
   38700: out<=1;
   38701: out<=1;
   38702: out<=1;
   38703: out<=1;
   38704: out<=0;
   38705: out<=0;
   38706: out<=1;
   38707: out<=1;
   38708: out<=1;
   38709: out<=0;
   38710: out<=1;
   38711: out<=0;
   38712: out<=1;
   38713: out<=0;
   38714: out<=0;
   38715: out<=1;
   38716: out<=0;
   38717: out<=0;
   38718: out<=0;
   38719: out<=0;
   38720: out<=1;
   38721: out<=1;
   38722: out<=0;
   38723: out<=0;
   38724: out<=0;
   38725: out<=1;
   38726: out<=0;
   38727: out<=1;
   38728: out<=0;
   38729: out<=1;
   38730: out<=1;
   38731: out<=0;
   38732: out<=1;
   38733: out<=1;
   38734: out<=1;
   38735: out<=1;
   38736: out<=1;
   38737: out<=1;
   38738: out<=0;
   38739: out<=0;
   38740: out<=0;
   38741: out<=1;
   38742: out<=0;
   38743: out<=1;
   38744: out<=0;
   38745: out<=1;
   38746: out<=1;
   38747: out<=0;
   38748: out<=1;
   38749: out<=1;
   38750: out<=1;
   38751: out<=1;
   38752: out<=0;
   38753: out<=0;
   38754: out<=1;
   38755: out<=1;
   38756: out<=1;
   38757: out<=0;
   38758: out<=1;
   38759: out<=0;
   38760: out<=1;
   38761: out<=0;
   38762: out<=0;
   38763: out<=1;
   38764: out<=0;
   38765: out<=0;
   38766: out<=0;
   38767: out<=0;
   38768: out<=0;
   38769: out<=0;
   38770: out<=1;
   38771: out<=1;
   38772: out<=1;
   38773: out<=0;
   38774: out<=1;
   38775: out<=0;
   38776: out<=1;
   38777: out<=0;
   38778: out<=0;
   38779: out<=1;
   38780: out<=0;
   38781: out<=0;
   38782: out<=0;
   38783: out<=0;
   38784: out<=0;
   38785: out<=0;
   38786: out<=1;
   38787: out<=1;
   38788: out<=1;
   38789: out<=0;
   38790: out<=1;
   38791: out<=0;
   38792: out<=1;
   38793: out<=0;
   38794: out<=0;
   38795: out<=1;
   38796: out<=0;
   38797: out<=0;
   38798: out<=0;
   38799: out<=0;
   38800: out<=0;
   38801: out<=0;
   38802: out<=1;
   38803: out<=1;
   38804: out<=1;
   38805: out<=0;
   38806: out<=1;
   38807: out<=0;
   38808: out<=1;
   38809: out<=0;
   38810: out<=0;
   38811: out<=1;
   38812: out<=0;
   38813: out<=0;
   38814: out<=0;
   38815: out<=0;
   38816: out<=0;
   38817: out<=0;
   38818: out<=1;
   38819: out<=1;
   38820: out<=1;
   38821: out<=0;
   38822: out<=1;
   38823: out<=0;
   38824: out<=1;
   38825: out<=0;
   38826: out<=0;
   38827: out<=1;
   38828: out<=0;
   38829: out<=0;
   38830: out<=0;
   38831: out<=0;
   38832: out<=0;
   38833: out<=0;
   38834: out<=1;
   38835: out<=1;
   38836: out<=1;
   38837: out<=0;
   38838: out<=1;
   38839: out<=0;
   38840: out<=1;
   38841: out<=0;
   38842: out<=0;
   38843: out<=1;
   38844: out<=0;
   38845: out<=0;
   38846: out<=0;
   38847: out<=0;
   38848: out<=0;
   38849: out<=0;
   38850: out<=1;
   38851: out<=1;
   38852: out<=1;
   38853: out<=0;
   38854: out<=1;
   38855: out<=0;
   38856: out<=1;
   38857: out<=0;
   38858: out<=0;
   38859: out<=1;
   38860: out<=0;
   38861: out<=0;
   38862: out<=0;
   38863: out<=0;
   38864: out<=1;
   38865: out<=1;
   38866: out<=0;
   38867: out<=0;
   38868: out<=0;
   38869: out<=1;
   38870: out<=0;
   38871: out<=1;
   38872: out<=0;
   38873: out<=1;
   38874: out<=1;
   38875: out<=0;
   38876: out<=1;
   38877: out<=1;
   38878: out<=1;
   38879: out<=1;
   38880: out<=1;
   38881: out<=1;
   38882: out<=0;
   38883: out<=0;
   38884: out<=0;
   38885: out<=1;
   38886: out<=0;
   38887: out<=1;
   38888: out<=0;
   38889: out<=1;
   38890: out<=1;
   38891: out<=0;
   38892: out<=1;
   38893: out<=1;
   38894: out<=1;
   38895: out<=1;
   38896: out<=0;
   38897: out<=0;
   38898: out<=1;
   38899: out<=1;
   38900: out<=1;
   38901: out<=0;
   38902: out<=1;
   38903: out<=0;
   38904: out<=1;
   38905: out<=0;
   38906: out<=0;
   38907: out<=1;
   38908: out<=0;
   38909: out<=0;
   38910: out<=0;
   38911: out<=0;
   38912: out<=1;
   38913: out<=1;
   38914: out<=0;
   38915: out<=0;
   38916: out<=0;
   38917: out<=1;
   38918: out<=0;
   38919: out<=1;
   38920: out<=1;
   38921: out<=0;
   38922: out<=0;
   38923: out<=1;
   38924: out<=0;
   38925: out<=0;
   38926: out<=0;
   38927: out<=0;
   38928: out<=0;
   38929: out<=0;
   38930: out<=1;
   38931: out<=1;
   38932: out<=1;
   38933: out<=0;
   38934: out<=1;
   38935: out<=0;
   38936: out<=0;
   38937: out<=1;
   38938: out<=1;
   38939: out<=0;
   38940: out<=1;
   38941: out<=1;
   38942: out<=1;
   38943: out<=1;
   38944: out<=0;
   38945: out<=0;
   38946: out<=1;
   38947: out<=1;
   38948: out<=1;
   38949: out<=0;
   38950: out<=1;
   38951: out<=0;
   38952: out<=0;
   38953: out<=1;
   38954: out<=1;
   38955: out<=0;
   38956: out<=1;
   38957: out<=1;
   38958: out<=1;
   38959: out<=1;
   38960: out<=1;
   38961: out<=1;
   38962: out<=0;
   38963: out<=0;
   38964: out<=0;
   38965: out<=1;
   38966: out<=0;
   38967: out<=1;
   38968: out<=1;
   38969: out<=0;
   38970: out<=0;
   38971: out<=1;
   38972: out<=0;
   38973: out<=0;
   38974: out<=0;
   38975: out<=0;
   38976: out<=1;
   38977: out<=1;
   38978: out<=0;
   38979: out<=0;
   38980: out<=0;
   38981: out<=1;
   38982: out<=0;
   38983: out<=1;
   38984: out<=1;
   38985: out<=0;
   38986: out<=0;
   38987: out<=1;
   38988: out<=0;
   38989: out<=0;
   38990: out<=0;
   38991: out<=0;
   38992: out<=1;
   38993: out<=1;
   38994: out<=0;
   38995: out<=0;
   38996: out<=0;
   38997: out<=1;
   38998: out<=0;
   38999: out<=1;
   39000: out<=1;
   39001: out<=0;
   39002: out<=0;
   39003: out<=1;
   39004: out<=0;
   39005: out<=0;
   39006: out<=0;
   39007: out<=0;
   39008: out<=1;
   39009: out<=1;
   39010: out<=0;
   39011: out<=0;
   39012: out<=0;
   39013: out<=1;
   39014: out<=0;
   39015: out<=1;
   39016: out<=1;
   39017: out<=0;
   39018: out<=0;
   39019: out<=1;
   39020: out<=0;
   39021: out<=0;
   39022: out<=0;
   39023: out<=0;
   39024: out<=1;
   39025: out<=1;
   39026: out<=0;
   39027: out<=0;
   39028: out<=0;
   39029: out<=1;
   39030: out<=0;
   39031: out<=1;
   39032: out<=1;
   39033: out<=0;
   39034: out<=0;
   39035: out<=1;
   39036: out<=0;
   39037: out<=0;
   39038: out<=0;
   39039: out<=0;
   39040: out<=0;
   39041: out<=0;
   39042: out<=1;
   39043: out<=1;
   39044: out<=1;
   39045: out<=0;
   39046: out<=1;
   39047: out<=0;
   39048: out<=0;
   39049: out<=1;
   39050: out<=1;
   39051: out<=0;
   39052: out<=1;
   39053: out<=1;
   39054: out<=1;
   39055: out<=1;
   39056: out<=0;
   39057: out<=0;
   39058: out<=1;
   39059: out<=1;
   39060: out<=1;
   39061: out<=0;
   39062: out<=1;
   39063: out<=0;
   39064: out<=0;
   39065: out<=1;
   39066: out<=1;
   39067: out<=0;
   39068: out<=1;
   39069: out<=1;
   39070: out<=1;
   39071: out<=1;
   39072: out<=1;
   39073: out<=1;
   39074: out<=0;
   39075: out<=0;
   39076: out<=0;
   39077: out<=1;
   39078: out<=0;
   39079: out<=1;
   39080: out<=1;
   39081: out<=0;
   39082: out<=0;
   39083: out<=1;
   39084: out<=0;
   39085: out<=0;
   39086: out<=0;
   39087: out<=0;
   39088: out<=1;
   39089: out<=1;
   39090: out<=0;
   39091: out<=0;
   39092: out<=0;
   39093: out<=1;
   39094: out<=0;
   39095: out<=1;
   39096: out<=1;
   39097: out<=0;
   39098: out<=0;
   39099: out<=1;
   39100: out<=0;
   39101: out<=0;
   39102: out<=0;
   39103: out<=0;
   39104: out<=0;
   39105: out<=0;
   39106: out<=1;
   39107: out<=1;
   39108: out<=1;
   39109: out<=0;
   39110: out<=1;
   39111: out<=0;
   39112: out<=0;
   39113: out<=1;
   39114: out<=1;
   39115: out<=0;
   39116: out<=1;
   39117: out<=1;
   39118: out<=1;
   39119: out<=1;
   39120: out<=1;
   39121: out<=1;
   39122: out<=0;
   39123: out<=0;
   39124: out<=0;
   39125: out<=1;
   39126: out<=0;
   39127: out<=1;
   39128: out<=1;
   39129: out<=0;
   39130: out<=0;
   39131: out<=1;
   39132: out<=0;
   39133: out<=0;
   39134: out<=0;
   39135: out<=0;
   39136: out<=0;
   39137: out<=0;
   39138: out<=1;
   39139: out<=1;
   39140: out<=1;
   39141: out<=0;
   39142: out<=1;
   39143: out<=0;
   39144: out<=0;
   39145: out<=1;
   39146: out<=1;
   39147: out<=0;
   39148: out<=1;
   39149: out<=1;
   39150: out<=1;
   39151: out<=1;
   39152: out<=1;
   39153: out<=1;
   39154: out<=0;
   39155: out<=0;
   39156: out<=0;
   39157: out<=1;
   39158: out<=0;
   39159: out<=1;
   39160: out<=1;
   39161: out<=0;
   39162: out<=0;
   39163: out<=1;
   39164: out<=0;
   39165: out<=0;
   39166: out<=0;
   39167: out<=0;
   39168: out<=0;
   39169: out<=1;
   39170: out<=0;
   39171: out<=1;
   39172: out<=0;
   39173: out<=0;
   39174: out<=1;
   39175: out<=1;
   39176: out<=1;
   39177: out<=1;
   39178: out<=1;
   39179: out<=1;
   39180: out<=1;
   39181: out<=0;
   39182: out<=0;
   39183: out<=1;
   39184: out<=0;
   39185: out<=1;
   39186: out<=0;
   39187: out<=1;
   39188: out<=0;
   39189: out<=0;
   39190: out<=1;
   39191: out<=1;
   39192: out<=1;
   39193: out<=1;
   39194: out<=1;
   39195: out<=1;
   39196: out<=1;
   39197: out<=0;
   39198: out<=0;
   39199: out<=1;
   39200: out<=0;
   39201: out<=1;
   39202: out<=0;
   39203: out<=1;
   39204: out<=0;
   39205: out<=0;
   39206: out<=1;
   39207: out<=1;
   39208: out<=1;
   39209: out<=1;
   39210: out<=1;
   39211: out<=1;
   39212: out<=1;
   39213: out<=0;
   39214: out<=0;
   39215: out<=1;
   39216: out<=0;
   39217: out<=1;
   39218: out<=0;
   39219: out<=1;
   39220: out<=0;
   39221: out<=0;
   39222: out<=1;
   39223: out<=1;
   39224: out<=1;
   39225: out<=1;
   39226: out<=1;
   39227: out<=1;
   39228: out<=1;
   39229: out<=0;
   39230: out<=0;
   39231: out<=1;
   39232: out<=0;
   39233: out<=1;
   39234: out<=0;
   39235: out<=1;
   39236: out<=0;
   39237: out<=0;
   39238: out<=1;
   39239: out<=1;
   39240: out<=1;
   39241: out<=1;
   39242: out<=1;
   39243: out<=1;
   39244: out<=1;
   39245: out<=0;
   39246: out<=0;
   39247: out<=1;
   39248: out<=1;
   39249: out<=0;
   39250: out<=1;
   39251: out<=0;
   39252: out<=1;
   39253: out<=1;
   39254: out<=0;
   39255: out<=0;
   39256: out<=0;
   39257: out<=0;
   39258: out<=0;
   39259: out<=0;
   39260: out<=0;
   39261: out<=1;
   39262: out<=1;
   39263: out<=0;
   39264: out<=1;
   39265: out<=0;
   39266: out<=1;
   39267: out<=0;
   39268: out<=1;
   39269: out<=1;
   39270: out<=0;
   39271: out<=0;
   39272: out<=0;
   39273: out<=0;
   39274: out<=0;
   39275: out<=0;
   39276: out<=0;
   39277: out<=1;
   39278: out<=1;
   39279: out<=0;
   39280: out<=0;
   39281: out<=1;
   39282: out<=0;
   39283: out<=1;
   39284: out<=0;
   39285: out<=0;
   39286: out<=1;
   39287: out<=1;
   39288: out<=1;
   39289: out<=1;
   39290: out<=1;
   39291: out<=1;
   39292: out<=1;
   39293: out<=0;
   39294: out<=0;
   39295: out<=1;
   39296: out<=1;
   39297: out<=0;
   39298: out<=1;
   39299: out<=0;
   39300: out<=1;
   39301: out<=1;
   39302: out<=0;
   39303: out<=0;
   39304: out<=0;
   39305: out<=0;
   39306: out<=0;
   39307: out<=0;
   39308: out<=0;
   39309: out<=1;
   39310: out<=1;
   39311: out<=0;
   39312: out<=0;
   39313: out<=1;
   39314: out<=0;
   39315: out<=1;
   39316: out<=0;
   39317: out<=0;
   39318: out<=1;
   39319: out<=1;
   39320: out<=1;
   39321: out<=1;
   39322: out<=1;
   39323: out<=1;
   39324: out<=1;
   39325: out<=0;
   39326: out<=0;
   39327: out<=1;
   39328: out<=1;
   39329: out<=0;
   39330: out<=1;
   39331: out<=0;
   39332: out<=1;
   39333: out<=1;
   39334: out<=0;
   39335: out<=0;
   39336: out<=0;
   39337: out<=0;
   39338: out<=0;
   39339: out<=0;
   39340: out<=0;
   39341: out<=1;
   39342: out<=1;
   39343: out<=0;
   39344: out<=0;
   39345: out<=1;
   39346: out<=0;
   39347: out<=1;
   39348: out<=0;
   39349: out<=0;
   39350: out<=1;
   39351: out<=1;
   39352: out<=1;
   39353: out<=1;
   39354: out<=1;
   39355: out<=1;
   39356: out<=1;
   39357: out<=0;
   39358: out<=0;
   39359: out<=1;
   39360: out<=1;
   39361: out<=0;
   39362: out<=1;
   39363: out<=0;
   39364: out<=1;
   39365: out<=1;
   39366: out<=0;
   39367: out<=0;
   39368: out<=0;
   39369: out<=0;
   39370: out<=0;
   39371: out<=0;
   39372: out<=0;
   39373: out<=1;
   39374: out<=1;
   39375: out<=0;
   39376: out<=1;
   39377: out<=0;
   39378: out<=1;
   39379: out<=0;
   39380: out<=1;
   39381: out<=1;
   39382: out<=0;
   39383: out<=0;
   39384: out<=0;
   39385: out<=0;
   39386: out<=0;
   39387: out<=0;
   39388: out<=0;
   39389: out<=1;
   39390: out<=1;
   39391: out<=0;
   39392: out<=0;
   39393: out<=1;
   39394: out<=0;
   39395: out<=1;
   39396: out<=0;
   39397: out<=0;
   39398: out<=1;
   39399: out<=1;
   39400: out<=1;
   39401: out<=1;
   39402: out<=1;
   39403: out<=1;
   39404: out<=1;
   39405: out<=0;
   39406: out<=0;
   39407: out<=1;
   39408: out<=0;
   39409: out<=1;
   39410: out<=0;
   39411: out<=1;
   39412: out<=0;
   39413: out<=0;
   39414: out<=1;
   39415: out<=1;
   39416: out<=1;
   39417: out<=1;
   39418: out<=1;
   39419: out<=1;
   39420: out<=1;
   39421: out<=0;
   39422: out<=0;
   39423: out<=1;
   39424: out<=1;
   39425: out<=0;
   39426: out<=0;
   39427: out<=1;
   39428: out<=1;
   39429: out<=1;
   39430: out<=1;
   39431: out<=1;
   39432: out<=1;
   39433: out<=1;
   39434: out<=0;
   39435: out<=0;
   39436: out<=1;
   39437: out<=0;
   39438: out<=1;
   39439: out<=0;
   39440: out<=1;
   39441: out<=0;
   39442: out<=0;
   39443: out<=1;
   39444: out<=1;
   39445: out<=1;
   39446: out<=1;
   39447: out<=1;
   39448: out<=1;
   39449: out<=1;
   39450: out<=0;
   39451: out<=0;
   39452: out<=1;
   39453: out<=0;
   39454: out<=1;
   39455: out<=0;
   39456: out<=0;
   39457: out<=1;
   39458: out<=1;
   39459: out<=0;
   39460: out<=0;
   39461: out<=0;
   39462: out<=0;
   39463: out<=0;
   39464: out<=0;
   39465: out<=0;
   39466: out<=1;
   39467: out<=1;
   39468: out<=0;
   39469: out<=1;
   39470: out<=0;
   39471: out<=1;
   39472: out<=0;
   39473: out<=1;
   39474: out<=1;
   39475: out<=0;
   39476: out<=0;
   39477: out<=0;
   39478: out<=0;
   39479: out<=0;
   39480: out<=0;
   39481: out<=0;
   39482: out<=1;
   39483: out<=1;
   39484: out<=0;
   39485: out<=1;
   39486: out<=0;
   39487: out<=1;
   39488: out<=1;
   39489: out<=0;
   39490: out<=0;
   39491: out<=1;
   39492: out<=1;
   39493: out<=1;
   39494: out<=1;
   39495: out<=1;
   39496: out<=1;
   39497: out<=1;
   39498: out<=0;
   39499: out<=0;
   39500: out<=1;
   39501: out<=0;
   39502: out<=1;
   39503: out<=0;
   39504: out<=0;
   39505: out<=1;
   39506: out<=1;
   39507: out<=0;
   39508: out<=0;
   39509: out<=0;
   39510: out<=0;
   39511: out<=0;
   39512: out<=0;
   39513: out<=0;
   39514: out<=1;
   39515: out<=1;
   39516: out<=0;
   39517: out<=1;
   39518: out<=0;
   39519: out<=1;
   39520: out<=1;
   39521: out<=0;
   39522: out<=0;
   39523: out<=1;
   39524: out<=1;
   39525: out<=1;
   39526: out<=1;
   39527: out<=1;
   39528: out<=1;
   39529: out<=1;
   39530: out<=0;
   39531: out<=0;
   39532: out<=1;
   39533: out<=0;
   39534: out<=1;
   39535: out<=0;
   39536: out<=0;
   39537: out<=1;
   39538: out<=1;
   39539: out<=0;
   39540: out<=0;
   39541: out<=0;
   39542: out<=0;
   39543: out<=0;
   39544: out<=0;
   39545: out<=0;
   39546: out<=1;
   39547: out<=1;
   39548: out<=0;
   39549: out<=1;
   39550: out<=0;
   39551: out<=1;
   39552: out<=0;
   39553: out<=1;
   39554: out<=1;
   39555: out<=0;
   39556: out<=0;
   39557: out<=0;
   39558: out<=0;
   39559: out<=0;
   39560: out<=0;
   39561: out<=0;
   39562: out<=1;
   39563: out<=1;
   39564: out<=0;
   39565: out<=1;
   39566: out<=0;
   39567: out<=1;
   39568: out<=1;
   39569: out<=0;
   39570: out<=0;
   39571: out<=1;
   39572: out<=1;
   39573: out<=1;
   39574: out<=1;
   39575: out<=1;
   39576: out<=1;
   39577: out<=1;
   39578: out<=0;
   39579: out<=0;
   39580: out<=1;
   39581: out<=0;
   39582: out<=1;
   39583: out<=0;
   39584: out<=1;
   39585: out<=0;
   39586: out<=0;
   39587: out<=1;
   39588: out<=1;
   39589: out<=1;
   39590: out<=1;
   39591: out<=1;
   39592: out<=1;
   39593: out<=1;
   39594: out<=0;
   39595: out<=0;
   39596: out<=1;
   39597: out<=0;
   39598: out<=1;
   39599: out<=0;
   39600: out<=0;
   39601: out<=1;
   39602: out<=1;
   39603: out<=0;
   39604: out<=0;
   39605: out<=0;
   39606: out<=0;
   39607: out<=0;
   39608: out<=0;
   39609: out<=0;
   39610: out<=1;
   39611: out<=1;
   39612: out<=0;
   39613: out<=1;
   39614: out<=0;
   39615: out<=1;
   39616: out<=0;
   39617: out<=1;
   39618: out<=1;
   39619: out<=0;
   39620: out<=0;
   39621: out<=0;
   39622: out<=0;
   39623: out<=0;
   39624: out<=0;
   39625: out<=0;
   39626: out<=1;
   39627: out<=1;
   39628: out<=0;
   39629: out<=1;
   39630: out<=0;
   39631: out<=1;
   39632: out<=0;
   39633: out<=1;
   39634: out<=1;
   39635: out<=0;
   39636: out<=0;
   39637: out<=0;
   39638: out<=0;
   39639: out<=0;
   39640: out<=0;
   39641: out<=0;
   39642: out<=1;
   39643: out<=1;
   39644: out<=0;
   39645: out<=1;
   39646: out<=0;
   39647: out<=1;
   39648: out<=0;
   39649: out<=1;
   39650: out<=1;
   39651: out<=0;
   39652: out<=0;
   39653: out<=0;
   39654: out<=0;
   39655: out<=0;
   39656: out<=0;
   39657: out<=0;
   39658: out<=1;
   39659: out<=1;
   39660: out<=0;
   39661: out<=1;
   39662: out<=0;
   39663: out<=1;
   39664: out<=0;
   39665: out<=1;
   39666: out<=1;
   39667: out<=0;
   39668: out<=0;
   39669: out<=0;
   39670: out<=0;
   39671: out<=0;
   39672: out<=0;
   39673: out<=0;
   39674: out<=1;
   39675: out<=1;
   39676: out<=0;
   39677: out<=1;
   39678: out<=0;
   39679: out<=1;
   39680: out<=0;
   39681: out<=0;
   39682: out<=0;
   39683: out<=0;
   39684: out<=1;
   39685: out<=0;
   39686: out<=0;
   39687: out<=1;
   39688: out<=1;
   39689: out<=0;
   39690: out<=1;
   39691: out<=0;
   39692: out<=0;
   39693: out<=0;
   39694: out<=1;
   39695: out<=1;
   39696: out<=1;
   39697: out<=1;
   39698: out<=1;
   39699: out<=1;
   39700: out<=0;
   39701: out<=1;
   39702: out<=1;
   39703: out<=0;
   39704: out<=0;
   39705: out<=1;
   39706: out<=0;
   39707: out<=1;
   39708: out<=1;
   39709: out<=1;
   39710: out<=0;
   39711: out<=0;
   39712: out<=0;
   39713: out<=0;
   39714: out<=0;
   39715: out<=0;
   39716: out<=1;
   39717: out<=0;
   39718: out<=0;
   39719: out<=1;
   39720: out<=1;
   39721: out<=0;
   39722: out<=1;
   39723: out<=0;
   39724: out<=0;
   39725: out<=0;
   39726: out<=1;
   39727: out<=1;
   39728: out<=1;
   39729: out<=1;
   39730: out<=1;
   39731: out<=1;
   39732: out<=0;
   39733: out<=1;
   39734: out<=1;
   39735: out<=0;
   39736: out<=0;
   39737: out<=1;
   39738: out<=0;
   39739: out<=1;
   39740: out<=1;
   39741: out<=1;
   39742: out<=0;
   39743: out<=0;
   39744: out<=0;
   39745: out<=0;
   39746: out<=0;
   39747: out<=0;
   39748: out<=1;
   39749: out<=0;
   39750: out<=0;
   39751: out<=1;
   39752: out<=1;
   39753: out<=0;
   39754: out<=1;
   39755: out<=0;
   39756: out<=0;
   39757: out<=0;
   39758: out<=1;
   39759: out<=1;
   39760: out<=0;
   39761: out<=0;
   39762: out<=0;
   39763: out<=0;
   39764: out<=1;
   39765: out<=0;
   39766: out<=0;
   39767: out<=1;
   39768: out<=1;
   39769: out<=0;
   39770: out<=1;
   39771: out<=0;
   39772: out<=0;
   39773: out<=0;
   39774: out<=1;
   39775: out<=1;
   39776: out<=1;
   39777: out<=1;
   39778: out<=1;
   39779: out<=1;
   39780: out<=0;
   39781: out<=1;
   39782: out<=1;
   39783: out<=0;
   39784: out<=0;
   39785: out<=1;
   39786: out<=0;
   39787: out<=1;
   39788: out<=1;
   39789: out<=1;
   39790: out<=0;
   39791: out<=0;
   39792: out<=1;
   39793: out<=1;
   39794: out<=1;
   39795: out<=1;
   39796: out<=0;
   39797: out<=1;
   39798: out<=1;
   39799: out<=0;
   39800: out<=0;
   39801: out<=1;
   39802: out<=0;
   39803: out<=1;
   39804: out<=1;
   39805: out<=1;
   39806: out<=0;
   39807: out<=0;
   39808: out<=1;
   39809: out<=1;
   39810: out<=1;
   39811: out<=1;
   39812: out<=0;
   39813: out<=1;
   39814: out<=1;
   39815: out<=0;
   39816: out<=0;
   39817: out<=1;
   39818: out<=0;
   39819: out<=1;
   39820: out<=1;
   39821: out<=1;
   39822: out<=0;
   39823: out<=0;
   39824: out<=1;
   39825: out<=1;
   39826: out<=1;
   39827: out<=1;
   39828: out<=0;
   39829: out<=1;
   39830: out<=1;
   39831: out<=0;
   39832: out<=0;
   39833: out<=1;
   39834: out<=0;
   39835: out<=1;
   39836: out<=1;
   39837: out<=1;
   39838: out<=0;
   39839: out<=0;
   39840: out<=1;
   39841: out<=1;
   39842: out<=1;
   39843: out<=1;
   39844: out<=0;
   39845: out<=1;
   39846: out<=1;
   39847: out<=0;
   39848: out<=0;
   39849: out<=1;
   39850: out<=0;
   39851: out<=1;
   39852: out<=1;
   39853: out<=1;
   39854: out<=0;
   39855: out<=0;
   39856: out<=1;
   39857: out<=1;
   39858: out<=1;
   39859: out<=1;
   39860: out<=0;
   39861: out<=1;
   39862: out<=1;
   39863: out<=0;
   39864: out<=0;
   39865: out<=1;
   39866: out<=0;
   39867: out<=1;
   39868: out<=1;
   39869: out<=1;
   39870: out<=0;
   39871: out<=0;
   39872: out<=1;
   39873: out<=1;
   39874: out<=1;
   39875: out<=1;
   39876: out<=0;
   39877: out<=1;
   39878: out<=1;
   39879: out<=0;
   39880: out<=0;
   39881: out<=1;
   39882: out<=0;
   39883: out<=1;
   39884: out<=1;
   39885: out<=1;
   39886: out<=0;
   39887: out<=0;
   39888: out<=0;
   39889: out<=0;
   39890: out<=0;
   39891: out<=0;
   39892: out<=1;
   39893: out<=0;
   39894: out<=0;
   39895: out<=1;
   39896: out<=1;
   39897: out<=0;
   39898: out<=1;
   39899: out<=0;
   39900: out<=0;
   39901: out<=0;
   39902: out<=1;
   39903: out<=1;
   39904: out<=0;
   39905: out<=0;
   39906: out<=0;
   39907: out<=0;
   39908: out<=1;
   39909: out<=0;
   39910: out<=0;
   39911: out<=1;
   39912: out<=1;
   39913: out<=0;
   39914: out<=1;
   39915: out<=0;
   39916: out<=0;
   39917: out<=0;
   39918: out<=1;
   39919: out<=1;
   39920: out<=1;
   39921: out<=1;
   39922: out<=1;
   39923: out<=1;
   39924: out<=0;
   39925: out<=1;
   39926: out<=1;
   39927: out<=0;
   39928: out<=0;
   39929: out<=1;
   39930: out<=0;
   39931: out<=1;
   39932: out<=1;
   39933: out<=1;
   39934: out<=0;
   39935: out<=0;
   39936: out<=1;
   39937: out<=0;
   39938: out<=1;
   39939: out<=0;
   39940: out<=0;
   39941: out<=0;
   39942: out<=1;
   39943: out<=1;
   39944: out<=1;
   39945: out<=1;
   39946: out<=1;
   39947: out<=1;
   39948: out<=0;
   39949: out<=1;
   39950: out<=1;
   39951: out<=0;
   39952: out<=0;
   39953: out<=1;
   39954: out<=0;
   39955: out<=1;
   39956: out<=1;
   39957: out<=1;
   39958: out<=0;
   39959: out<=0;
   39960: out<=0;
   39961: out<=0;
   39962: out<=0;
   39963: out<=0;
   39964: out<=1;
   39965: out<=0;
   39966: out<=0;
   39967: out<=1;
   39968: out<=0;
   39969: out<=1;
   39970: out<=0;
   39971: out<=1;
   39972: out<=1;
   39973: out<=1;
   39974: out<=0;
   39975: out<=0;
   39976: out<=0;
   39977: out<=0;
   39978: out<=0;
   39979: out<=0;
   39980: out<=1;
   39981: out<=0;
   39982: out<=0;
   39983: out<=1;
   39984: out<=1;
   39985: out<=0;
   39986: out<=1;
   39987: out<=0;
   39988: out<=0;
   39989: out<=0;
   39990: out<=1;
   39991: out<=1;
   39992: out<=1;
   39993: out<=1;
   39994: out<=1;
   39995: out<=1;
   39996: out<=0;
   39997: out<=1;
   39998: out<=1;
   39999: out<=0;
   40000: out<=1;
   40001: out<=0;
   40002: out<=1;
   40003: out<=0;
   40004: out<=0;
   40005: out<=0;
   40006: out<=1;
   40007: out<=1;
   40008: out<=1;
   40009: out<=1;
   40010: out<=1;
   40011: out<=1;
   40012: out<=0;
   40013: out<=1;
   40014: out<=1;
   40015: out<=0;
   40016: out<=1;
   40017: out<=0;
   40018: out<=1;
   40019: out<=0;
   40020: out<=0;
   40021: out<=0;
   40022: out<=1;
   40023: out<=1;
   40024: out<=1;
   40025: out<=1;
   40026: out<=1;
   40027: out<=1;
   40028: out<=0;
   40029: out<=1;
   40030: out<=1;
   40031: out<=0;
   40032: out<=1;
   40033: out<=0;
   40034: out<=1;
   40035: out<=0;
   40036: out<=0;
   40037: out<=0;
   40038: out<=1;
   40039: out<=1;
   40040: out<=1;
   40041: out<=1;
   40042: out<=1;
   40043: out<=1;
   40044: out<=0;
   40045: out<=1;
   40046: out<=1;
   40047: out<=0;
   40048: out<=1;
   40049: out<=0;
   40050: out<=1;
   40051: out<=0;
   40052: out<=0;
   40053: out<=0;
   40054: out<=1;
   40055: out<=1;
   40056: out<=1;
   40057: out<=1;
   40058: out<=1;
   40059: out<=1;
   40060: out<=0;
   40061: out<=1;
   40062: out<=1;
   40063: out<=0;
   40064: out<=0;
   40065: out<=1;
   40066: out<=0;
   40067: out<=1;
   40068: out<=1;
   40069: out<=1;
   40070: out<=0;
   40071: out<=0;
   40072: out<=0;
   40073: out<=0;
   40074: out<=0;
   40075: out<=0;
   40076: out<=1;
   40077: out<=0;
   40078: out<=0;
   40079: out<=1;
   40080: out<=0;
   40081: out<=1;
   40082: out<=0;
   40083: out<=1;
   40084: out<=1;
   40085: out<=1;
   40086: out<=0;
   40087: out<=0;
   40088: out<=0;
   40089: out<=0;
   40090: out<=0;
   40091: out<=0;
   40092: out<=1;
   40093: out<=0;
   40094: out<=0;
   40095: out<=1;
   40096: out<=1;
   40097: out<=0;
   40098: out<=1;
   40099: out<=0;
   40100: out<=0;
   40101: out<=0;
   40102: out<=1;
   40103: out<=1;
   40104: out<=1;
   40105: out<=1;
   40106: out<=1;
   40107: out<=1;
   40108: out<=0;
   40109: out<=1;
   40110: out<=1;
   40111: out<=0;
   40112: out<=1;
   40113: out<=0;
   40114: out<=1;
   40115: out<=0;
   40116: out<=0;
   40117: out<=0;
   40118: out<=1;
   40119: out<=1;
   40120: out<=1;
   40121: out<=1;
   40122: out<=1;
   40123: out<=1;
   40124: out<=0;
   40125: out<=1;
   40126: out<=1;
   40127: out<=0;
   40128: out<=0;
   40129: out<=1;
   40130: out<=0;
   40131: out<=1;
   40132: out<=1;
   40133: out<=1;
   40134: out<=0;
   40135: out<=0;
   40136: out<=0;
   40137: out<=0;
   40138: out<=0;
   40139: out<=0;
   40140: out<=1;
   40141: out<=0;
   40142: out<=0;
   40143: out<=1;
   40144: out<=1;
   40145: out<=0;
   40146: out<=1;
   40147: out<=0;
   40148: out<=0;
   40149: out<=0;
   40150: out<=1;
   40151: out<=1;
   40152: out<=1;
   40153: out<=1;
   40154: out<=1;
   40155: out<=1;
   40156: out<=0;
   40157: out<=1;
   40158: out<=1;
   40159: out<=0;
   40160: out<=0;
   40161: out<=1;
   40162: out<=0;
   40163: out<=1;
   40164: out<=1;
   40165: out<=1;
   40166: out<=0;
   40167: out<=0;
   40168: out<=0;
   40169: out<=0;
   40170: out<=0;
   40171: out<=0;
   40172: out<=1;
   40173: out<=0;
   40174: out<=0;
   40175: out<=1;
   40176: out<=1;
   40177: out<=0;
   40178: out<=1;
   40179: out<=0;
   40180: out<=0;
   40181: out<=0;
   40182: out<=1;
   40183: out<=1;
   40184: out<=1;
   40185: out<=1;
   40186: out<=1;
   40187: out<=1;
   40188: out<=0;
   40189: out<=1;
   40190: out<=1;
   40191: out<=0;
   40192: out<=1;
   40193: out<=1;
   40194: out<=0;
   40195: out<=0;
   40196: out<=1;
   40197: out<=0;
   40198: out<=1;
   40199: out<=0;
   40200: out<=0;
   40201: out<=1;
   40202: out<=1;
   40203: out<=0;
   40204: out<=0;
   40205: out<=0;
   40206: out<=0;
   40207: out<=0;
   40208: out<=1;
   40209: out<=1;
   40210: out<=0;
   40211: out<=0;
   40212: out<=1;
   40213: out<=0;
   40214: out<=1;
   40215: out<=0;
   40216: out<=0;
   40217: out<=1;
   40218: out<=1;
   40219: out<=0;
   40220: out<=0;
   40221: out<=0;
   40222: out<=0;
   40223: out<=0;
   40224: out<=1;
   40225: out<=1;
   40226: out<=0;
   40227: out<=0;
   40228: out<=1;
   40229: out<=0;
   40230: out<=1;
   40231: out<=0;
   40232: out<=0;
   40233: out<=1;
   40234: out<=1;
   40235: out<=0;
   40236: out<=0;
   40237: out<=0;
   40238: out<=0;
   40239: out<=0;
   40240: out<=1;
   40241: out<=1;
   40242: out<=0;
   40243: out<=0;
   40244: out<=1;
   40245: out<=0;
   40246: out<=1;
   40247: out<=0;
   40248: out<=0;
   40249: out<=1;
   40250: out<=1;
   40251: out<=0;
   40252: out<=0;
   40253: out<=0;
   40254: out<=0;
   40255: out<=0;
   40256: out<=1;
   40257: out<=1;
   40258: out<=0;
   40259: out<=0;
   40260: out<=1;
   40261: out<=0;
   40262: out<=1;
   40263: out<=0;
   40264: out<=0;
   40265: out<=1;
   40266: out<=1;
   40267: out<=0;
   40268: out<=0;
   40269: out<=0;
   40270: out<=0;
   40271: out<=0;
   40272: out<=0;
   40273: out<=0;
   40274: out<=1;
   40275: out<=1;
   40276: out<=0;
   40277: out<=1;
   40278: out<=0;
   40279: out<=1;
   40280: out<=1;
   40281: out<=0;
   40282: out<=0;
   40283: out<=1;
   40284: out<=1;
   40285: out<=1;
   40286: out<=1;
   40287: out<=1;
   40288: out<=0;
   40289: out<=0;
   40290: out<=1;
   40291: out<=1;
   40292: out<=0;
   40293: out<=1;
   40294: out<=0;
   40295: out<=1;
   40296: out<=1;
   40297: out<=0;
   40298: out<=0;
   40299: out<=1;
   40300: out<=1;
   40301: out<=1;
   40302: out<=1;
   40303: out<=1;
   40304: out<=1;
   40305: out<=1;
   40306: out<=0;
   40307: out<=0;
   40308: out<=1;
   40309: out<=0;
   40310: out<=1;
   40311: out<=0;
   40312: out<=0;
   40313: out<=1;
   40314: out<=1;
   40315: out<=0;
   40316: out<=0;
   40317: out<=0;
   40318: out<=0;
   40319: out<=0;
   40320: out<=0;
   40321: out<=0;
   40322: out<=1;
   40323: out<=1;
   40324: out<=0;
   40325: out<=1;
   40326: out<=0;
   40327: out<=1;
   40328: out<=1;
   40329: out<=0;
   40330: out<=0;
   40331: out<=1;
   40332: out<=1;
   40333: out<=1;
   40334: out<=1;
   40335: out<=1;
   40336: out<=1;
   40337: out<=1;
   40338: out<=0;
   40339: out<=0;
   40340: out<=1;
   40341: out<=0;
   40342: out<=1;
   40343: out<=0;
   40344: out<=0;
   40345: out<=1;
   40346: out<=1;
   40347: out<=0;
   40348: out<=0;
   40349: out<=0;
   40350: out<=0;
   40351: out<=0;
   40352: out<=0;
   40353: out<=0;
   40354: out<=1;
   40355: out<=1;
   40356: out<=0;
   40357: out<=1;
   40358: out<=0;
   40359: out<=1;
   40360: out<=1;
   40361: out<=0;
   40362: out<=0;
   40363: out<=1;
   40364: out<=1;
   40365: out<=1;
   40366: out<=1;
   40367: out<=1;
   40368: out<=1;
   40369: out<=1;
   40370: out<=0;
   40371: out<=0;
   40372: out<=1;
   40373: out<=0;
   40374: out<=1;
   40375: out<=0;
   40376: out<=0;
   40377: out<=1;
   40378: out<=1;
   40379: out<=0;
   40380: out<=0;
   40381: out<=0;
   40382: out<=0;
   40383: out<=0;
   40384: out<=0;
   40385: out<=0;
   40386: out<=1;
   40387: out<=1;
   40388: out<=0;
   40389: out<=1;
   40390: out<=0;
   40391: out<=1;
   40392: out<=1;
   40393: out<=0;
   40394: out<=0;
   40395: out<=1;
   40396: out<=1;
   40397: out<=1;
   40398: out<=1;
   40399: out<=1;
   40400: out<=0;
   40401: out<=0;
   40402: out<=1;
   40403: out<=1;
   40404: out<=0;
   40405: out<=1;
   40406: out<=0;
   40407: out<=1;
   40408: out<=1;
   40409: out<=0;
   40410: out<=0;
   40411: out<=1;
   40412: out<=1;
   40413: out<=1;
   40414: out<=1;
   40415: out<=1;
   40416: out<=1;
   40417: out<=1;
   40418: out<=0;
   40419: out<=0;
   40420: out<=1;
   40421: out<=0;
   40422: out<=1;
   40423: out<=0;
   40424: out<=0;
   40425: out<=1;
   40426: out<=1;
   40427: out<=0;
   40428: out<=0;
   40429: out<=0;
   40430: out<=0;
   40431: out<=0;
   40432: out<=1;
   40433: out<=1;
   40434: out<=0;
   40435: out<=0;
   40436: out<=1;
   40437: out<=0;
   40438: out<=1;
   40439: out<=0;
   40440: out<=0;
   40441: out<=1;
   40442: out<=1;
   40443: out<=0;
   40444: out<=0;
   40445: out<=0;
   40446: out<=0;
   40447: out<=0;
   40448: out<=0;
   40449: out<=0;
   40450: out<=0;
   40451: out<=0;
   40452: out<=0;
   40453: out<=1;
   40454: out<=1;
   40455: out<=0;
   40456: out<=0;
   40457: out<=1;
   40458: out<=0;
   40459: out<=1;
   40460: out<=0;
   40461: out<=0;
   40462: out<=1;
   40463: out<=1;
   40464: out<=0;
   40465: out<=0;
   40466: out<=0;
   40467: out<=0;
   40468: out<=0;
   40469: out<=1;
   40470: out<=1;
   40471: out<=0;
   40472: out<=0;
   40473: out<=1;
   40474: out<=0;
   40475: out<=1;
   40476: out<=0;
   40477: out<=0;
   40478: out<=1;
   40479: out<=1;
   40480: out<=1;
   40481: out<=1;
   40482: out<=1;
   40483: out<=1;
   40484: out<=1;
   40485: out<=0;
   40486: out<=0;
   40487: out<=1;
   40488: out<=1;
   40489: out<=0;
   40490: out<=1;
   40491: out<=0;
   40492: out<=1;
   40493: out<=1;
   40494: out<=0;
   40495: out<=0;
   40496: out<=1;
   40497: out<=1;
   40498: out<=1;
   40499: out<=1;
   40500: out<=1;
   40501: out<=0;
   40502: out<=0;
   40503: out<=1;
   40504: out<=1;
   40505: out<=0;
   40506: out<=1;
   40507: out<=0;
   40508: out<=1;
   40509: out<=1;
   40510: out<=0;
   40511: out<=0;
   40512: out<=0;
   40513: out<=0;
   40514: out<=0;
   40515: out<=0;
   40516: out<=0;
   40517: out<=1;
   40518: out<=1;
   40519: out<=0;
   40520: out<=0;
   40521: out<=1;
   40522: out<=0;
   40523: out<=1;
   40524: out<=0;
   40525: out<=0;
   40526: out<=1;
   40527: out<=1;
   40528: out<=1;
   40529: out<=1;
   40530: out<=1;
   40531: out<=1;
   40532: out<=1;
   40533: out<=0;
   40534: out<=0;
   40535: out<=1;
   40536: out<=1;
   40537: out<=0;
   40538: out<=1;
   40539: out<=0;
   40540: out<=1;
   40541: out<=1;
   40542: out<=0;
   40543: out<=0;
   40544: out<=0;
   40545: out<=0;
   40546: out<=0;
   40547: out<=0;
   40548: out<=0;
   40549: out<=1;
   40550: out<=1;
   40551: out<=0;
   40552: out<=0;
   40553: out<=1;
   40554: out<=0;
   40555: out<=1;
   40556: out<=0;
   40557: out<=0;
   40558: out<=1;
   40559: out<=1;
   40560: out<=1;
   40561: out<=1;
   40562: out<=1;
   40563: out<=1;
   40564: out<=1;
   40565: out<=0;
   40566: out<=0;
   40567: out<=1;
   40568: out<=1;
   40569: out<=0;
   40570: out<=1;
   40571: out<=0;
   40572: out<=1;
   40573: out<=1;
   40574: out<=0;
   40575: out<=0;
   40576: out<=1;
   40577: out<=1;
   40578: out<=1;
   40579: out<=1;
   40580: out<=1;
   40581: out<=0;
   40582: out<=0;
   40583: out<=1;
   40584: out<=1;
   40585: out<=0;
   40586: out<=1;
   40587: out<=0;
   40588: out<=1;
   40589: out<=1;
   40590: out<=0;
   40591: out<=0;
   40592: out<=0;
   40593: out<=0;
   40594: out<=0;
   40595: out<=0;
   40596: out<=0;
   40597: out<=1;
   40598: out<=1;
   40599: out<=0;
   40600: out<=0;
   40601: out<=1;
   40602: out<=0;
   40603: out<=1;
   40604: out<=0;
   40605: out<=0;
   40606: out<=1;
   40607: out<=1;
   40608: out<=0;
   40609: out<=0;
   40610: out<=0;
   40611: out<=0;
   40612: out<=0;
   40613: out<=1;
   40614: out<=1;
   40615: out<=0;
   40616: out<=0;
   40617: out<=1;
   40618: out<=0;
   40619: out<=1;
   40620: out<=0;
   40621: out<=0;
   40622: out<=1;
   40623: out<=1;
   40624: out<=1;
   40625: out<=1;
   40626: out<=1;
   40627: out<=1;
   40628: out<=1;
   40629: out<=0;
   40630: out<=0;
   40631: out<=1;
   40632: out<=1;
   40633: out<=0;
   40634: out<=1;
   40635: out<=0;
   40636: out<=1;
   40637: out<=1;
   40638: out<=0;
   40639: out<=0;
   40640: out<=1;
   40641: out<=1;
   40642: out<=1;
   40643: out<=1;
   40644: out<=1;
   40645: out<=0;
   40646: out<=0;
   40647: out<=1;
   40648: out<=1;
   40649: out<=0;
   40650: out<=1;
   40651: out<=0;
   40652: out<=1;
   40653: out<=1;
   40654: out<=0;
   40655: out<=0;
   40656: out<=1;
   40657: out<=1;
   40658: out<=1;
   40659: out<=1;
   40660: out<=1;
   40661: out<=0;
   40662: out<=0;
   40663: out<=1;
   40664: out<=1;
   40665: out<=0;
   40666: out<=1;
   40667: out<=0;
   40668: out<=1;
   40669: out<=1;
   40670: out<=0;
   40671: out<=0;
   40672: out<=1;
   40673: out<=1;
   40674: out<=1;
   40675: out<=1;
   40676: out<=1;
   40677: out<=0;
   40678: out<=0;
   40679: out<=1;
   40680: out<=1;
   40681: out<=0;
   40682: out<=1;
   40683: out<=0;
   40684: out<=1;
   40685: out<=1;
   40686: out<=0;
   40687: out<=0;
   40688: out<=1;
   40689: out<=1;
   40690: out<=1;
   40691: out<=1;
   40692: out<=1;
   40693: out<=0;
   40694: out<=0;
   40695: out<=1;
   40696: out<=1;
   40697: out<=0;
   40698: out<=1;
   40699: out<=0;
   40700: out<=1;
   40701: out<=1;
   40702: out<=0;
   40703: out<=0;
   40704: out<=0;
   40705: out<=1;
   40706: out<=1;
   40707: out<=0;
   40708: out<=1;
   40709: out<=1;
   40710: out<=1;
   40711: out<=1;
   40712: out<=1;
   40713: out<=1;
   40714: out<=0;
   40715: out<=0;
   40716: out<=0;
   40717: out<=1;
   40718: out<=0;
   40719: out<=1;
   40720: out<=1;
   40721: out<=0;
   40722: out<=0;
   40723: out<=1;
   40724: out<=0;
   40725: out<=0;
   40726: out<=0;
   40727: out<=0;
   40728: out<=0;
   40729: out<=0;
   40730: out<=1;
   40731: out<=1;
   40732: out<=1;
   40733: out<=0;
   40734: out<=1;
   40735: out<=0;
   40736: out<=0;
   40737: out<=1;
   40738: out<=1;
   40739: out<=0;
   40740: out<=1;
   40741: out<=1;
   40742: out<=1;
   40743: out<=1;
   40744: out<=1;
   40745: out<=1;
   40746: out<=0;
   40747: out<=0;
   40748: out<=0;
   40749: out<=1;
   40750: out<=0;
   40751: out<=1;
   40752: out<=1;
   40753: out<=0;
   40754: out<=0;
   40755: out<=1;
   40756: out<=0;
   40757: out<=0;
   40758: out<=0;
   40759: out<=0;
   40760: out<=0;
   40761: out<=0;
   40762: out<=1;
   40763: out<=1;
   40764: out<=1;
   40765: out<=0;
   40766: out<=1;
   40767: out<=0;
   40768: out<=0;
   40769: out<=1;
   40770: out<=1;
   40771: out<=0;
   40772: out<=1;
   40773: out<=1;
   40774: out<=1;
   40775: out<=1;
   40776: out<=1;
   40777: out<=1;
   40778: out<=0;
   40779: out<=0;
   40780: out<=0;
   40781: out<=1;
   40782: out<=0;
   40783: out<=1;
   40784: out<=0;
   40785: out<=1;
   40786: out<=1;
   40787: out<=0;
   40788: out<=1;
   40789: out<=1;
   40790: out<=1;
   40791: out<=1;
   40792: out<=1;
   40793: out<=1;
   40794: out<=0;
   40795: out<=0;
   40796: out<=0;
   40797: out<=1;
   40798: out<=0;
   40799: out<=1;
   40800: out<=1;
   40801: out<=0;
   40802: out<=0;
   40803: out<=1;
   40804: out<=0;
   40805: out<=0;
   40806: out<=0;
   40807: out<=0;
   40808: out<=0;
   40809: out<=0;
   40810: out<=1;
   40811: out<=1;
   40812: out<=1;
   40813: out<=0;
   40814: out<=1;
   40815: out<=0;
   40816: out<=1;
   40817: out<=0;
   40818: out<=0;
   40819: out<=1;
   40820: out<=0;
   40821: out<=0;
   40822: out<=0;
   40823: out<=0;
   40824: out<=0;
   40825: out<=0;
   40826: out<=1;
   40827: out<=1;
   40828: out<=1;
   40829: out<=0;
   40830: out<=1;
   40831: out<=0;
   40832: out<=1;
   40833: out<=0;
   40834: out<=0;
   40835: out<=1;
   40836: out<=0;
   40837: out<=0;
   40838: out<=0;
   40839: out<=0;
   40840: out<=0;
   40841: out<=0;
   40842: out<=1;
   40843: out<=1;
   40844: out<=1;
   40845: out<=0;
   40846: out<=1;
   40847: out<=0;
   40848: out<=1;
   40849: out<=0;
   40850: out<=0;
   40851: out<=1;
   40852: out<=0;
   40853: out<=0;
   40854: out<=0;
   40855: out<=0;
   40856: out<=0;
   40857: out<=0;
   40858: out<=1;
   40859: out<=1;
   40860: out<=1;
   40861: out<=0;
   40862: out<=1;
   40863: out<=0;
   40864: out<=1;
   40865: out<=0;
   40866: out<=0;
   40867: out<=1;
   40868: out<=0;
   40869: out<=0;
   40870: out<=0;
   40871: out<=0;
   40872: out<=0;
   40873: out<=0;
   40874: out<=1;
   40875: out<=1;
   40876: out<=1;
   40877: out<=0;
   40878: out<=1;
   40879: out<=0;
   40880: out<=1;
   40881: out<=0;
   40882: out<=0;
   40883: out<=1;
   40884: out<=0;
   40885: out<=0;
   40886: out<=0;
   40887: out<=0;
   40888: out<=0;
   40889: out<=0;
   40890: out<=1;
   40891: out<=1;
   40892: out<=1;
   40893: out<=0;
   40894: out<=1;
   40895: out<=0;
   40896: out<=1;
   40897: out<=0;
   40898: out<=0;
   40899: out<=1;
   40900: out<=0;
   40901: out<=0;
   40902: out<=0;
   40903: out<=0;
   40904: out<=0;
   40905: out<=0;
   40906: out<=1;
   40907: out<=1;
   40908: out<=1;
   40909: out<=0;
   40910: out<=1;
   40911: out<=0;
   40912: out<=0;
   40913: out<=1;
   40914: out<=1;
   40915: out<=0;
   40916: out<=1;
   40917: out<=1;
   40918: out<=1;
   40919: out<=1;
   40920: out<=1;
   40921: out<=1;
   40922: out<=0;
   40923: out<=0;
   40924: out<=0;
   40925: out<=1;
   40926: out<=0;
   40927: out<=1;
   40928: out<=0;
   40929: out<=1;
   40930: out<=1;
   40931: out<=0;
   40932: out<=1;
   40933: out<=1;
   40934: out<=1;
   40935: out<=1;
   40936: out<=1;
   40937: out<=1;
   40938: out<=0;
   40939: out<=0;
   40940: out<=0;
   40941: out<=1;
   40942: out<=0;
   40943: out<=1;
   40944: out<=1;
   40945: out<=0;
   40946: out<=0;
   40947: out<=1;
   40948: out<=0;
   40949: out<=0;
   40950: out<=0;
   40951: out<=0;
   40952: out<=0;
   40953: out<=0;
   40954: out<=1;
   40955: out<=1;
   40956: out<=1;
   40957: out<=0;
   40958: out<=1;
   40959: out<=0;
   40960: out<=0;
   40961: out<=1;
   40962: out<=0;
   40963: out<=1;
   40964: out<=1;
   40965: out<=1;
   40966: out<=0;
   40967: out<=0;
   40968: out<=0;
   40969: out<=0;
   40970: out<=0;
   40971: out<=0;
   40972: out<=1;
   40973: out<=0;
   40974: out<=0;
   40975: out<=1;
   40976: out<=1;
   40977: out<=0;
   40978: out<=1;
   40979: out<=0;
   40980: out<=0;
   40981: out<=0;
   40982: out<=1;
   40983: out<=1;
   40984: out<=1;
   40985: out<=1;
   40986: out<=1;
   40987: out<=1;
   40988: out<=0;
   40989: out<=1;
   40990: out<=1;
   40991: out<=0;
   40992: out<=0;
   40993: out<=1;
   40994: out<=0;
   40995: out<=1;
   40996: out<=1;
   40997: out<=1;
   40998: out<=0;
   40999: out<=0;
   41000: out<=0;
   41001: out<=0;
   41002: out<=0;
   41003: out<=0;
   41004: out<=1;
   41005: out<=0;
   41006: out<=0;
   41007: out<=1;
   41008: out<=1;
   41009: out<=0;
   41010: out<=1;
   41011: out<=0;
   41012: out<=0;
   41013: out<=0;
   41014: out<=1;
   41015: out<=1;
   41016: out<=1;
   41017: out<=1;
   41018: out<=1;
   41019: out<=1;
   41020: out<=0;
   41021: out<=1;
   41022: out<=1;
   41023: out<=0;
   41024: out<=0;
   41025: out<=1;
   41026: out<=0;
   41027: out<=1;
   41028: out<=1;
   41029: out<=1;
   41030: out<=0;
   41031: out<=0;
   41032: out<=0;
   41033: out<=0;
   41034: out<=0;
   41035: out<=0;
   41036: out<=1;
   41037: out<=0;
   41038: out<=0;
   41039: out<=1;
   41040: out<=0;
   41041: out<=1;
   41042: out<=0;
   41043: out<=1;
   41044: out<=1;
   41045: out<=1;
   41046: out<=0;
   41047: out<=0;
   41048: out<=0;
   41049: out<=0;
   41050: out<=0;
   41051: out<=0;
   41052: out<=1;
   41053: out<=0;
   41054: out<=0;
   41055: out<=1;
   41056: out<=1;
   41057: out<=0;
   41058: out<=1;
   41059: out<=0;
   41060: out<=0;
   41061: out<=0;
   41062: out<=1;
   41063: out<=1;
   41064: out<=1;
   41065: out<=1;
   41066: out<=1;
   41067: out<=1;
   41068: out<=0;
   41069: out<=1;
   41070: out<=1;
   41071: out<=0;
   41072: out<=1;
   41073: out<=0;
   41074: out<=1;
   41075: out<=0;
   41076: out<=0;
   41077: out<=0;
   41078: out<=1;
   41079: out<=1;
   41080: out<=1;
   41081: out<=1;
   41082: out<=1;
   41083: out<=1;
   41084: out<=0;
   41085: out<=1;
   41086: out<=1;
   41087: out<=0;
   41088: out<=0;
   41089: out<=1;
   41090: out<=0;
   41091: out<=1;
   41092: out<=1;
   41093: out<=1;
   41094: out<=0;
   41095: out<=0;
   41096: out<=0;
   41097: out<=0;
   41098: out<=0;
   41099: out<=0;
   41100: out<=1;
   41101: out<=0;
   41102: out<=0;
   41103: out<=1;
   41104: out<=0;
   41105: out<=1;
   41106: out<=0;
   41107: out<=1;
   41108: out<=1;
   41109: out<=1;
   41110: out<=0;
   41111: out<=0;
   41112: out<=0;
   41113: out<=0;
   41114: out<=0;
   41115: out<=0;
   41116: out<=1;
   41117: out<=0;
   41118: out<=0;
   41119: out<=1;
   41120: out<=0;
   41121: out<=1;
   41122: out<=0;
   41123: out<=1;
   41124: out<=1;
   41125: out<=1;
   41126: out<=0;
   41127: out<=0;
   41128: out<=0;
   41129: out<=0;
   41130: out<=0;
   41131: out<=0;
   41132: out<=1;
   41133: out<=0;
   41134: out<=0;
   41135: out<=1;
   41136: out<=0;
   41137: out<=1;
   41138: out<=0;
   41139: out<=1;
   41140: out<=1;
   41141: out<=1;
   41142: out<=0;
   41143: out<=0;
   41144: out<=0;
   41145: out<=0;
   41146: out<=0;
   41147: out<=0;
   41148: out<=1;
   41149: out<=0;
   41150: out<=0;
   41151: out<=1;
   41152: out<=0;
   41153: out<=1;
   41154: out<=0;
   41155: out<=1;
   41156: out<=1;
   41157: out<=1;
   41158: out<=0;
   41159: out<=0;
   41160: out<=0;
   41161: out<=0;
   41162: out<=0;
   41163: out<=0;
   41164: out<=1;
   41165: out<=0;
   41166: out<=0;
   41167: out<=1;
   41168: out<=1;
   41169: out<=0;
   41170: out<=1;
   41171: out<=0;
   41172: out<=0;
   41173: out<=0;
   41174: out<=1;
   41175: out<=1;
   41176: out<=1;
   41177: out<=1;
   41178: out<=1;
   41179: out<=1;
   41180: out<=0;
   41181: out<=1;
   41182: out<=1;
   41183: out<=0;
   41184: out<=1;
   41185: out<=0;
   41186: out<=1;
   41187: out<=0;
   41188: out<=0;
   41189: out<=0;
   41190: out<=1;
   41191: out<=1;
   41192: out<=1;
   41193: out<=1;
   41194: out<=1;
   41195: out<=1;
   41196: out<=0;
   41197: out<=1;
   41198: out<=1;
   41199: out<=0;
   41200: out<=0;
   41201: out<=1;
   41202: out<=0;
   41203: out<=1;
   41204: out<=1;
   41205: out<=1;
   41206: out<=0;
   41207: out<=0;
   41208: out<=0;
   41209: out<=0;
   41210: out<=0;
   41211: out<=0;
   41212: out<=1;
   41213: out<=0;
   41214: out<=0;
   41215: out<=1;
   41216: out<=0;
   41217: out<=0;
   41218: out<=1;
   41219: out<=1;
   41220: out<=0;
   41221: out<=1;
   41222: out<=0;
   41223: out<=1;
   41224: out<=1;
   41225: out<=0;
   41226: out<=0;
   41227: out<=1;
   41228: out<=1;
   41229: out<=1;
   41230: out<=1;
   41231: out<=1;
   41232: out<=0;
   41233: out<=0;
   41234: out<=1;
   41235: out<=1;
   41236: out<=0;
   41237: out<=1;
   41238: out<=0;
   41239: out<=1;
   41240: out<=1;
   41241: out<=0;
   41242: out<=0;
   41243: out<=1;
   41244: out<=1;
   41245: out<=1;
   41246: out<=1;
   41247: out<=1;
   41248: out<=1;
   41249: out<=1;
   41250: out<=0;
   41251: out<=0;
   41252: out<=1;
   41253: out<=0;
   41254: out<=1;
   41255: out<=0;
   41256: out<=0;
   41257: out<=1;
   41258: out<=1;
   41259: out<=0;
   41260: out<=0;
   41261: out<=0;
   41262: out<=0;
   41263: out<=0;
   41264: out<=1;
   41265: out<=1;
   41266: out<=0;
   41267: out<=0;
   41268: out<=1;
   41269: out<=0;
   41270: out<=1;
   41271: out<=0;
   41272: out<=0;
   41273: out<=1;
   41274: out<=1;
   41275: out<=0;
   41276: out<=0;
   41277: out<=0;
   41278: out<=0;
   41279: out<=0;
   41280: out<=0;
   41281: out<=0;
   41282: out<=1;
   41283: out<=1;
   41284: out<=0;
   41285: out<=1;
   41286: out<=0;
   41287: out<=1;
   41288: out<=1;
   41289: out<=0;
   41290: out<=0;
   41291: out<=1;
   41292: out<=1;
   41293: out<=1;
   41294: out<=1;
   41295: out<=1;
   41296: out<=1;
   41297: out<=1;
   41298: out<=0;
   41299: out<=0;
   41300: out<=1;
   41301: out<=0;
   41302: out<=1;
   41303: out<=0;
   41304: out<=0;
   41305: out<=1;
   41306: out<=1;
   41307: out<=0;
   41308: out<=0;
   41309: out<=0;
   41310: out<=0;
   41311: out<=0;
   41312: out<=0;
   41313: out<=0;
   41314: out<=1;
   41315: out<=1;
   41316: out<=0;
   41317: out<=1;
   41318: out<=0;
   41319: out<=1;
   41320: out<=1;
   41321: out<=0;
   41322: out<=0;
   41323: out<=1;
   41324: out<=1;
   41325: out<=1;
   41326: out<=1;
   41327: out<=1;
   41328: out<=1;
   41329: out<=1;
   41330: out<=0;
   41331: out<=0;
   41332: out<=1;
   41333: out<=0;
   41334: out<=1;
   41335: out<=0;
   41336: out<=0;
   41337: out<=1;
   41338: out<=1;
   41339: out<=0;
   41340: out<=0;
   41341: out<=0;
   41342: out<=0;
   41343: out<=0;
   41344: out<=0;
   41345: out<=0;
   41346: out<=1;
   41347: out<=1;
   41348: out<=0;
   41349: out<=1;
   41350: out<=0;
   41351: out<=1;
   41352: out<=1;
   41353: out<=0;
   41354: out<=0;
   41355: out<=1;
   41356: out<=1;
   41357: out<=1;
   41358: out<=1;
   41359: out<=1;
   41360: out<=1;
   41361: out<=1;
   41362: out<=0;
   41363: out<=0;
   41364: out<=1;
   41365: out<=0;
   41366: out<=1;
   41367: out<=0;
   41368: out<=0;
   41369: out<=1;
   41370: out<=1;
   41371: out<=0;
   41372: out<=0;
   41373: out<=0;
   41374: out<=0;
   41375: out<=0;
   41376: out<=1;
   41377: out<=1;
   41378: out<=0;
   41379: out<=0;
   41380: out<=1;
   41381: out<=0;
   41382: out<=1;
   41383: out<=0;
   41384: out<=0;
   41385: out<=1;
   41386: out<=1;
   41387: out<=0;
   41388: out<=0;
   41389: out<=0;
   41390: out<=0;
   41391: out<=0;
   41392: out<=0;
   41393: out<=0;
   41394: out<=1;
   41395: out<=1;
   41396: out<=0;
   41397: out<=1;
   41398: out<=0;
   41399: out<=1;
   41400: out<=1;
   41401: out<=0;
   41402: out<=0;
   41403: out<=1;
   41404: out<=1;
   41405: out<=1;
   41406: out<=1;
   41407: out<=1;
   41408: out<=0;
   41409: out<=0;
   41410: out<=1;
   41411: out<=1;
   41412: out<=0;
   41413: out<=1;
   41414: out<=0;
   41415: out<=1;
   41416: out<=1;
   41417: out<=0;
   41418: out<=0;
   41419: out<=1;
   41420: out<=1;
   41421: out<=1;
   41422: out<=1;
   41423: out<=1;
   41424: out<=0;
   41425: out<=0;
   41426: out<=1;
   41427: out<=1;
   41428: out<=0;
   41429: out<=1;
   41430: out<=0;
   41431: out<=1;
   41432: out<=1;
   41433: out<=0;
   41434: out<=0;
   41435: out<=1;
   41436: out<=1;
   41437: out<=1;
   41438: out<=1;
   41439: out<=1;
   41440: out<=0;
   41441: out<=0;
   41442: out<=1;
   41443: out<=1;
   41444: out<=0;
   41445: out<=1;
   41446: out<=0;
   41447: out<=1;
   41448: out<=1;
   41449: out<=0;
   41450: out<=0;
   41451: out<=1;
   41452: out<=1;
   41453: out<=1;
   41454: out<=1;
   41455: out<=1;
   41456: out<=0;
   41457: out<=0;
   41458: out<=1;
   41459: out<=1;
   41460: out<=0;
   41461: out<=1;
   41462: out<=0;
   41463: out<=1;
   41464: out<=1;
   41465: out<=0;
   41466: out<=0;
   41467: out<=1;
   41468: out<=1;
   41469: out<=1;
   41470: out<=1;
   41471: out<=1;
   41472: out<=0;
   41473: out<=0;
   41474: out<=0;
   41475: out<=0;
   41476: out<=0;
   41477: out<=1;
   41478: out<=1;
   41479: out<=0;
   41480: out<=0;
   41481: out<=1;
   41482: out<=0;
   41483: out<=1;
   41484: out<=0;
   41485: out<=0;
   41486: out<=1;
   41487: out<=1;
   41488: out<=0;
   41489: out<=0;
   41490: out<=0;
   41491: out<=0;
   41492: out<=0;
   41493: out<=1;
   41494: out<=1;
   41495: out<=0;
   41496: out<=0;
   41497: out<=1;
   41498: out<=0;
   41499: out<=1;
   41500: out<=0;
   41501: out<=0;
   41502: out<=1;
   41503: out<=1;
   41504: out<=0;
   41505: out<=0;
   41506: out<=0;
   41507: out<=0;
   41508: out<=0;
   41509: out<=1;
   41510: out<=1;
   41511: out<=0;
   41512: out<=0;
   41513: out<=1;
   41514: out<=0;
   41515: out<=1;
   41516: out<=0;
   41517: out<=0;
   41518: out<=1;
   41519: out<=1;
   41520: out<=0;
   41521: out<=0;
   41522: out<=0;
   41523: out<=0;
   41524: out<=0;
   41525: out<=1;
   41526: out<=1;
   41527: out<=0;
   41528: out<=0;
   41529: out<=1;
   41530: out<=0;
   41531: out<=1;
   41532: out<=0;
   41533: out<=0;
   41534: out<=1;
   41535: out<=1;
   41536: out<=0;
   41537: out<=0;
   41538: out<=0;
   41539: out<=0;
   41540: out<=0;
   41541: out<=1;
   41542: out<=1;
   41543: out<=0;
   41544: out<=0;
   41545: out<=1;
   41546: out<=0;
   41547: out<=1;
   41548: out<=0;
   41549: out<=0;
   41550: out<=1;
   41551: out<=1;
   41552: out<=1;
   41553: out<=1;
   41554: out<=1;
   41555: out<=1;
   41556: out<=1;
   41557: out<=0;
   41558: out<=0;
   41559: out<=1;
   41560: out<=1;
   41561: out<=0;
   41562: out<=1;
   41563: out<=0;
   41564: out<=1;
   41565: out<=1;
   41566: out<=0;
   41567: out<=0;
   41568: out<=1;
   41569: out<=1;
   41570: out<=1;
   41571: out<=1;
   41572: out<=1;
   41573: out<=0;
   41574: out<=0;
   41575: out<=1;
   41576: out<=1;
   41577: out<=0;
   41578: out<=1;
   41579: out<=0;
   41580: out<=1;
   41581: out<=1;
   41582: out<=0;
   41583: out<=0;
   41584: out<=0;
   41585: out<=0;
   41586: out<=0;
   41587: out<=0;
   41588: out<=0;
   41589: out<=1;
   41590: out<=1;
   41591: out<=0;
   41592: out<=0;
   41593: out<=1;
   41594: out<=0;
   41595: out<=1;
   41596: out<=0;
   41597: out<=0;
   41598: out<=1;
   41599: out<=1;
   41600: out<=0;
   41601: out<=0;
   41602: out<=0;
   41603: out<=0;
   41604: out<=0;
   41605: out<=1;
   41606: out<=1;
   41607: out<=0;
   41608: out<=0;
   41609: out<=1;
   41610: out<=0;
   41611: out<=1;
   41612: out<=0;
   41613: out<=0;
   41614: out<=1;
   41615: out<=1;
   41616: out<=1;
   41617: out<=1;
   41618: out<=1;
   41619: out<=1;
   41620: out<=1;
   41621: out<=0;
   41622: out<=0;
   41623: out<=1;
   41624: out<=1;
   41625: out<=0;
   41626: out<=1;
   41627: out<=0;
   41628: out<=1;
   41629: out<=1;
   41630: out<=0;
   41631: out<=0;
   41632: out<=0;
   41633: out<=0;
   41634: out<=0;
   41635: out<=0;
   41636: out<=0;
   41637: out<=1;
   41638: out<=1;
   41639: out<=0;
   41640: out<=0;
   41641: out<=1;
   41642: out<=0;
   41643: out<=1;
   41644: out<=0;
   41645: out<=0;
   41646: out<=1;
   41647: out<=1;
   41648: out<=1;
   41649: out<=1;
   41650: out<=1;
   41651: out<=1;
   41652: out<=1;
   41653: out<=0;
   41654: out<=0;
   41655: out<=1;
   41656: out<=1;
   41657: out<=0;
   41658: out<=1;
   41659: out<=0;
   41660: out<=1;
   41661: out<=1;
   41662: out<=0;
   41663: out<=0;
   41664: out<=0;
   41665: out<=0;
   41666: out<=0;
   41667: out<=0;
   41668: out<=0;
   41669: out<=1;
   41670: out<=1;
   41671: out<=0;
   41672: out<=0;
   41673: out<=1;
   41674: out<=0;
   41675: out<=1;
   41676: out<=0;
   41677: out<=0;
   41678: out<=1;
   41679: out<=1;
   41680: out<=0;
   41681: out<=0;
   41682: out<=0;
   41683: out<=0;
   41684: out<=0;
   41685: out<=1;
   41686: out<=1;
   41687: out<=0;
   41688: out<=0;
   41689: out<=1;
   41690: out<=0;
   41691: out<=1;
   41692: out<=0;
   41693: out<=0;
   41694: out<=1;
   41695: out<=1;
   41696: out<=1;
   41697: out<=1;
   41698: out<=1;
   41699: out<=1;
   41700: out<=1;
   41701: out<=0;
   41702: out<=0;
   41703: out<=1;
   41704: out<=1;
   41705: out<=0;
   41706: out<=1;
   41707: out<=0;
   41708: out<=1;
   41709: out<=1;
   41710: out<=0;
   41711: out<=0;
   41712: out<=1;
   41713: out<=1;
   41714: out<=1;
   41715: out<=1;
   41716: out<=1;
   41717: out<=0;
   41718: out<=0;
   41719: out<=1;
   41720: out<=1;
   41721: out<=0;
   41722: out<=1;
   41723: out<=0;
   41724: out<=1;
   41725: out<=1;
   41726: out<=0;
   41727: out<=0;
   41728: out<=0;
   41729: out<=1;
   41730: out<=1;
   41731: out<=0;
   41732: out<=1;
   41733: out<=1;
   41734: out<=1;
   41735: out<=1;
   41736: out<=1;
   41737: out<=1;
   41738: out<=0;
   41739: out<=0;
   41740: out<=0;
   41741: out<=1;
   41742: out<=0;
   41743: out<=1;
   41744: out<=1;
   41745: out<=0;
   41746: out<=0;
   41747: out<=1;
   41748: out<=0;
   41749: out<=0;
   41750: out<=0;
   41751: out<=0;
   41752: out<=0;
   41753: out<=0;
   41754: out<=1;
   41755: out<=1;
   41756: out<=1;
   41757: out<=0;
   41758: out<=1;
   41759: out<=0;
   41760: out<=1;
   41761: out<=0;
   41762: out<=0;
   41763: out<=1;
   41764: out<=0;
   41765: out<=0;
   41766: out<=0;
   41767: out<=0;
   41768: out<=0;
   41769: out<=0;
   41770: out<=1;
   41771: out<=1;
   41772: out<=1;
   41773: out<=0;
   41774: out<=1;
   41775: out<=0;
   41776: out<=0;
   41777: out<=1;
   41778: out<=1;
   41779: out<=0;
   41780: out<=1;
   41781: out<=1;
   41782: out<=1;
   41783: out<=1;
   41784: out<=1;
   41785: out<=1;
   41786: out<=0;
   41787: out<=0;
   41788: out<=0;
   41789: out<=1;
   41790: out<=0;
   41791: out<=1;
   41792: out<=0;
   41793: out<=1;
   41794: out<=1;
   41795: out<=0;
   41796: out<=1;
   41797: out<=1;
   41798: out<=1;
   41799: out<=1;
   41800: out<=1;
   41801: out<=1;
   41802: out<=0;
   41803: out<=0;
   41804: out<=0;
   41805: out<=1;
   41806: out<=0;
   41807: out<=1;
   41808: out<=0;
   41809: out<=1;
   41810: out<=1;
   41811: out<=0;
   41812: out<=1;
   41813: out<=1;
   41814: out<=1;
   41815: out<=1;
   41816: out<=1;
   41817: out<=1;
   41818: out<=0;
   41819: out<=0;
   41820: out<=0;
   41821: out<=1;
   41822: out<=0;
   41823: out<=1;
   41824: out<=0;
   41825: out<=1;
   41826: out<=1;
   41827: out<=0;
   41828: out<=1;
   41829: out<=1;
   41830: out<=1;
   41831: out<=1;
   41832: out<=1;
   41833: out<=1;
   41834: out<=0;
   41835: out<=0;
   41836: out<=0;
   41837: out<=1;
   41838: out<=0;
   41839: out<=1;
   41840: out<=0;
   41841: out<=1;
   41842: out<=1;
   41843: out<=0;
   41844: out<=1;
   41845: out<=1;
   41846: out<=1;
   41847: out<=1;
   41848: out<=1;
   41849: out<=1;
   41850: out<=0;
   41851: out<=0;
   41852: out<=0;
   41853: out<=1;
   41854: out<=0;
   41855: out<=1;
   41856: out<=0;
   41857: out<=1;
   41858: out<=1;
   41859: out<=0;
   41860: out<=1;
   41861: out<=1;
   41862: out<=1;
   41863: out<=1;
   41864: out<=1;
   41865: out<=1;
   41866: out<=0;
   41867: out<=0;
   41868: out<=0;
   41869: out<=1;
   41870: out<=0;
   41871: out<=1;
   41872: out<=0;
   41873: out<=1;
   41874: out<=1;
   41875: out<=0;
   41876: out<=1;
   41877: out<=1;
   41878: out<=1;
   41879: out<=1;
   41880: out<=1;
   41881: out<=1;
   41882: out<=0;
   41883: out<=0;
   41884: out<=0;
   41885: out<=1;
   41886: out<=0;
   41887: out<=1;
   41888: out<=1;
   41889: out<=0;
   41890: out<=0;
   41891: out<=1;
   41892: out<=0;
   41893: out<=0;
   41894: out<=0;
   41895: out<=0;
   41896: out<=0;
   41897: out<=0;
   41898: out<=1;
   41899: out<=1;
   41900: out<=1;
   41901: out<=0;
   41902: out<=1;
   41903: out<=0;
   41904: out<=1;
   41905: out<=0;
   41906: out<=0;
   41907: out<=1;
   41908: out<=0;
   41909: out<=0;
   41910: out<=0;
   41911: out<=0;
   41912: out<=0;
   41913: out<=0;
   41914: out<=1;
   41915: out<=1;
   41916: out<=1;
   41917: out<=0;
   41918: out<=1;
   41919: out<=0;
   41920: out<=0;
   41921: out<=1;
   41922: out<=1;
   41923: out<=0;
   41924: out<=1;
   41925: out<=1;
   41926: out<=1;
   41927: out<=1;
   41928: out<=1;
   41929: out<=1;
   41930: out<=0;
   41931: out<=0;
   41932: out<=0;
   41933: out<=1;
   41934: out<=0;
   41935: out<=1;
   41936: out<=1;
   41937: out<=0;
   41938: out<=0;
   41939: out<=1;
   41940: out<=0;
   41941: out<=0;
   41942: out<=0;
   41943: out<=0;
   41944: out<=0;
   41945: out<=0;
   41946: out<=1;
   41947: out<=1;
   41948: out<=1;
   41949: out<=0;
   41950: out<=1;
   41951: out<=0;
   41952: out<=0;
   41953: out<=1;
   41954: out<=1;
   41955: out<=0;
   41956: out<=1;
   41957: out<=1;
   41958: out<=1;
   41959: out<=1;
   41960: out<=1;
   41961: out<=1;
   41962: out<=0;
   41963: out<=0;
   41964: out<=0;
   41965: out<=1;
   41966: out<=0;
   41967: out<=1;
   41968: out<=1;
   41969: out<=0;
   41970: out<=0;
   41971: out<=1;
   41972: out<=0;
   41973: out<=0;
   41974: out<=0;
   41975: out<=0;
   41976: out<=0;
   41977: out<=0;
   41978: out<=1;
   41979: out<=1;
   41980: out<=1;
   41981: out<=0;
   41982: out<=1;
   41983: out<=0;
   41984: out<=0;
   41985: out<=0;
   41986: out<=1;
   41987: out<=1;
   41988: out<=1;
   41989: out<=0;
   41990: out<=1;
   41991: out<=0;
   41992: out<=0;
   41993: out<=1;
   41994: out<=1;
   41995: out<=0;
   41996: out<=1;
   41997: out<=1;
   41998: out<=1;
   41999: out<=1;
   42000: out<=1;
   42001: out<=1;
   42002: out<=0;
   42003: out<=0;
   42004: out<=0;
   42005: out<=1;
   42006: out<=0;
   42007: out<=1;
   42008: out<=1;
   42009: out<=0;
   42010: out<=0;
   42011: out<=1;
   42012: out<=0;
   42013: out<=0;
   42014: out<=0;
   42015: out<=0;
   42016: out<=0;
   42017: out<=0;
   42018: out<=1;
   42019: out<=1;
   42020: out<=1;
   42021: out<=0;
   42022: out<=1;
   42023: out<=0;
   42024: out<=0;
   42025: out<=1;
   42026: out<=1;
   42027: out<=0;
   42028: out<=1;
   42029: out<=1;
   42030: out<=1;
   42031: out<=1;
   42032: out<=1;
   42033: out<=1;
   42034: out<=0;
   42035: out<=0;
   42036: out<=0;
   42037: out<=1;
   42038: out<=0;
   42039: out<=1;
   42040: out<=1;
   42041: out<=0;
   42042: out<=0;
   42043: out<=1;
   42044: out<=0;
   42045: out<=0;
   42046: out<=0;
   42047: out<=0;
   42048: out<=0;
   42049: out<=0;
   42050: out<=1;
   42051: out<=1;
   42052: out<=1;
   42053: out<=0;
   42054: out<=1;
   42055: out<=0;
   42056: out<=0;
   42057: out<=1;
   42058: out<=1;
   42059: out<=0;
   42060: out<=1;
   42061: out<=1;
   42062: out<=1;
   42063: out<=1;
   42064: out<=0;
   42065: out<=0;
   42066: out<=1;
   42067: out<=1;
   42068: out<=1;
   42069: out<=0;
   42070: out<=1;
   42071: out<=0;
   42072: out<=0;
   42073: out<=1;
   42074: out<=1;
   42075: out<=0;
   42076: out<=1;
   42077: out<=1;
   42078: out<=1;
   42079: out<=1;
   42080: out<=1;
   42081: out<=1;
   42082: out<=0;
   42083: out<=0;
   42084: out<=0;
   42085: out<=1;
   42086: out<=0;
   42087: out<=1;
   42088: out<=1;
   42089: out<=0;
   42090: out<=0;
   42091: out<=1;
   42092: out<=0;
   42093: out<=0;
   42094: out<=0;
   42095: out<=0;
   42096: out<=1;
   42097: out<=1;
   42098: out<=0;
   42099: out<=0;
   42100: out<=0;
   42101: out<=1;
   42102: out<=0;
   42103: out<=1;
   42104: out<=1;
   42105: out<=0;
   42106: out<=0;
   42107: out<=1;
   42108: out<=0;
   42109: out<=0;
   42110: out<=0;
   42111: out<=0;
   42112: out<=0;
   42113: out<=0;
   42114: out<=1;
   42115: out<=1;
   42116: out<=1;
   42117: out<=0;
   42118: out<=1;
   42119: out<=0;
   42120: out<=0;
   42121: out<=1;
   42122: out<=1;
   42123: out<=0;
   42124: out<=1;
   42125: out<=1;
   42126: out<=1;
   42127: out<=1;
   42128: out<=0;
   42129: out<=0;
   42130: out<=1;
   42131: out<=1;
   42132: out<=1;
   42133: out<=0;
   42134: out<=1;
   42135: out<=0;
   42136: out<=0;
   42137: out<=1;
   42138: out<=1;
   42139: out<=0;
   42140: out<=1;
   42141: out<=1;
   42142: out<=1;
   42143: out<=1;
   42144: out<=0;
   42145: out<=0;
   42146: out<=1;
   42147: out<=1;
   42148: out<=1;
   42149: out<=0;
   42150: out<=1;
   42151: out<=0;
   42152: out<=0;
   42153: out<=1;
   42154: out<=1;
   42155: out<=0;
   42156: out<=1;
   42157: out<=1;
   42158: out<=1;
   42159: out<=1;
   42160: out<=0;
   42161: out<=0;
   42162: out<=1;
   42163: out<=1;
   42164: out<=1;
   42165: out<=0;
   42166: out<=1;
   42167: out<=0;
   42168: out<=0;
   42169: out<=1;
   42170: out<=1;
   42171: out<=0;
   42172: out<=1;
   42173: out<=1;
   42174: out<=1;
   42175: out<=1;
   42176: out<=0;
   42177: out<=0;
   42178: out<=1;
   42179: out<=1;
   42180: out<=1;
   42181: out<=0;
   42182: out<=1;
   42183: out<=0;
   42184: out<=0;
   42185: out<=1;
   42186: out<=1;
   42187: out<=0;
   42188: out<=1;
   42189: out<=1;
   42190: out<=1;
   42191: out<=1;
   42192: out<=1;
   42193: out<=1;
   42194: out<=0;
   42195: out<=0;
   42196: out<=0;
   42197: out<=1;
   42198: out<=0;
   42199: out<=1;
   42200: out<=1;
   42201: out<=0;
   42202: out<=0;
   42203: out<=1;
   42204: out<=0;
   42205: out<=0;
   42206: out<=0;
   42207: out<=0;
   42208: out<=1;
   42209: out<=1;
   42210: out<=0;
   42211: out<=0;
   42212: out<=0;
   42213: out<=1;
   42214: out<=0;
   42215: out<=1;
   42216: out<=1;
   42217: out<=0;
   42218: out<=0;
   42219: out<=1;
   42220: out<=0;
   42221: out<=0;
   42222: out<=0;
   42223: out<=0;
   42224: out<=0;
   42225: out<=0;
   42226: out<=1;
   42227: out<=1;
   42228: out<=1;
   42229: out<=0;
   42230: out<=1;
   42231: out<=0;
   42232: out<=0;
   42233: out<=1;
   42234: out<=1;
   42235: out<=0;
   42236: out<=1;
   42237: out<=1;
   42238: out<=1;
   42239: out<=1;
   42240: out<=1;
   42241: out<=0;
   42242: out<=1;
   42243: out<=0;
   42244: out<=1;
   42245: out<=1;
   42246: out<=0;
   42247: out<=0;
   42248: out<=0;
   42249: out<=0;
   42250: out<=0;
   42251: out<=0;
   42252: out<=0;
   42253: out<=1;
   42254: out<=1;
   42255: out<=0;
   42256: out<=1;
   42257: out<=0;
   42258: out<=1;
   42259: out<=0;
   42260: out<=1;
   42261: out<=1;
   42262: out<=0;
   42263: out<=0;
   42264: out<=0;
   42265: out<=0;
   42266: out<=0;
   42267: out<=0;
   42268: out<=0;
   42269: out<=1;
   42270: out<=1;
   42271: out<=0;
   42272: out<=0;
   42273: out<=1;
   42274: out<=0;
   42275: out<=1;
   42276: out<=0;
   42277: out<=0;
   42278: out<=1;
   42279: out<=1;
   42280: out<=1;
   42281: out<=1;
   42282: out<=1;
   42283: out<=1;
   42284: out<=1;
   42285: out<=0;
   42286: out<=0;
   42287: out<=1;
   42288: out<=0;
   42289: out<=1;
   42290: out<=0;
   42291: out<=1;
   42292: out<=0;
   42293: out<=0;
   42294: out<=1;
   42295: out<=1;
   42296: out<=1;
   42297: out<=1;
   42298: out<=1;
   42299: out<=1;
   42300: out<=1;
   42301: out<=0;
   42302: out<=0;
   42303: out<=1;
   42304: out<=1;
   42305: out<=0;
   42306: out<=1;
   42307: out<=0;
   42308: out<=1;
   42309: out<=1;
   42310: out<=0;
   42311: out<=0;
   42312: out<=0;
   42313: out<=0;
   42314: out<=0;
   42315: out<=0;
   42316: out<=0;
   42317: out<=1;
   42318: out<=1;
   42319: out<=0;
   42320: out<=0;
   42321: out<=1;
   42322: out<=0;
   42323: out<=1;
   42324: out<=0;
   42325: out<=0;
   42326: out<=1;
   42327: out<=1;
   42328: out<=1;
   42329: out<=1;
   42330: out<=1;
   42331: out<=1;
   42332: out<=1;
   42333: out<=0;
   42334: out<=0;
   42335: out<=1;
   42336: out<=1;
   42337: out<=0;
   42338: out<=1;
   42339: out<=0;
   42340: out<=1;
   42341: out<=1;
   42342: out<=0;
   42343: out<=0;
   42344: out<=0;
   42345: out<=0;
   42346: out<=0;
   42347: out<=0;
   42348: out<=0;
   42349: out<=1;
   42350: out<=1;
   42351: out<=0;
   42352: out<=0;
   42353: out<=1;
   42354: out<=0;
   42355: out<=1;
   42356: out<=0;
   42357: out<=0;
   42358: out<=1;
   42359: out<=1;
   42360: out<=1;
   42361: out<=1;
   42362: out<=1;
   42363: out<=1;
   42364: out<=1;
   42365: out<=0;
   42366: out<=0;
   42367: out<=1;
   42368: out<=1;
   42369: out<=0;
   42370: out<=1;
   42371: out<=0;
   42372: out<=1;
   42373: out<=1;
   42374: out<=0;
   42375: out<=0;
   42376: out<=0;
   42377: out<=0;
   42378: out<=0;
   42379: out<=0;
   42380: out<=0;
   42381: out<=1;
   42382: out<=1;
   42383: out<=0;
   42384: out<=0;
   42385: out<=1;
   42386: out<=0;
   42387: out<=1;
   42388: out<=0;
   42389: out<=0;
   42390: out<=1;
   42391: out<=1;
   42392: out<=1;
   42393: out<=1;
   42394: out<=1;
   42395: out<=1;
   42396: out<=1;
   42397: out<=0;
   42398: out<=0;
   42399: out<=1;
   42400: out<=0;
   42401: out<=1;
   42402: out<=0;
   42403: out<=1;
   42404: out<=0;
   42405: out<=0;
   42406: out<=1;
   42407: out<=1;
   42408: out<=1;
   42409: out<=1;
   42410: out<=1;
   42411: out<=1;
   42412: out<=1;
   42413: out<=0;
   42414: out<=0;
   42415: out<=1;
   42416: out<=1;
   42417: out<=0;
   42418: out<=1;
   42419: out<=0;
   42420: out<=1;
   42421: out<=1;
   42422: out<=0;
   42423: out<=0;
   42424: out<=0;
   42425: out<=0;
   42426: out<=0;
   42427: out<=0;
   42428: out<=0;
   42429: out<=1;
   42430: out<=1;
   42431: out<=0;
   42432: out<=1;
   42433: out<=0;
   42434: out<=1;
   42435: out<=0;
   42436: out<=1;
   42437: out<=1;
   42438: out<=0;
   42439: out<=0;
   42440: out<=0;
   42441: out<=0;
   42442: out<=0;
   42443: out<=0;
   42444: out<=0;
   42445: out<=1;
   42446: out<=1;
   42447: out<=0;
   42448: out<=1;
   42449: out<=0;
   42450: out<=1;
   42451: out<=0;
   42452: out<=1;
   42453: out<=1;
   42454: out<=0;
   42455: out<=0;
   42456: out<=0;
   42457: out<=0;
   42458: out<=0;
   42459: out<=0;
   42460: out<=0;
   42461: out<=1;
   42462: out<=1;
   42463: out<=0;
   42464: out<=1;
   42465: out<=0;
   42466: out<=1;
   42467: out<=0;
   42468: out<=1;
   42469: out<=1;
   42470: out<=0;
   42471: out<=0;
   42472: out<=0;
   42473: out<=0;
   42474: out<=0;
   42475: out<=0;
   42476: out<=0;
   42477: out<=1;
   42478: out<=1;
   42479: out<=0;
   42480: out<=1;
   42481: out<=0;
   42482: out<=1;
   42483: out<=0;
   42484: out<=1;
   42485: out<=1;
   42486: out<=0;
   42487: out<=0;
   42488: out<=0;
   42489: out<=0;
   42490: out<=0;
   42491: out<=0;
   42492: out<=0;
   42493: out<=1;
   42494: out<=1;
   42495: out<=0;
   42496: out<=1;
   42497: out<=0;
   42498: out<=0;
   42499: out<=1;
   42500: out<=1;
   42501: out<=1;
   42502: out<=1;
   42503: out<=1;
   42504: out<=1;
   42505: out<=1;
   42506: out<=0;
   42507: out<=0;
   42508: out<=1;
   42509: out<=0;
   42510: out<=1;
   42511: out<=0;
   42512: out<=1;
   42513: out<=0;
   42514: out<=0;
   42515: out<=1;
   42516: out<=1;
   42517: out<=1;
   42518: out<=1;
   42519: out<=1;
   42520: out<=1;
   42521: out<=1;
   42522: out<=0;
   42523: out<=0;
   42524: out<=1;
   42525: out<=0;
   42526: out<=1;
   42527: out<=0;
   42528: out<=1;
   42529: out<=0;
   42530: out<=0;
   42531: out<=1;
   42532: out<=1;
   42533: out<=1;
   42534: out<=1;
   42535: out<=1;
   42536: out<=1;
   42537: out<=1;
   42538: out<=0;
   42539: out<=0;
   42540: out<=1;
   42541: out<=0;
   42542: out<=1;
   42543: out<=0;
   42544: out<=1;
   42545: out<=0;
   42546: out<=0;
   42547: out<=1;
   42548: out<=1;
   42549: out<=1;
   42550: out<=1;
   42551: out<=1;
   42552: out<=1;
   42553: out<=1;
   42554: out<=0;
   42555: out<=0;
   42556: out<=1;
   42557: out<=0;
   42558: out<=1;
   42559: out<=0;
   42560: out<=1;
   42561: out<=0;
   42562: out<=0;
   42563: out<=1;
   42564: out<=1;
   42565: out<=1;
   42566: out<=1;
   42567: out<=1;
   42568: out<=1;
   42569: out<=1;
   42570: out<=0;
   42571: out<=0;
   42572: out<=1;
   42573: out<=0;
   42574: out<=1;
   42575: out<=0;
   42576: out<=0;
   42577: out<=1;
   42578: out<=1;
   42579: out<=0;
   42580: out<=0;
   42581: out<=0;
   42582: out<=0;
   42583: out<=0;
   42584: out<=0;
   42585: out<=0;
   42586: out<=1;
   42587: out<=1;
   42588: out<=0;
   42589: out<=1;
   42590: out<=0;
   42591: out<=1;
   42592: out<=0;
   42593: out<=1;
   42594: out<=1;
   42595: out<=0;
   42596: out<=0;
   42597: out<=0;
   42598: out<=0;
   42599: out<=0;
   42600: out<=0;
   42601: out<=0;
   42602: out<=1;
   42603: out<=1;
   42604: out<=0;
   42605: out<=1;
   42606: out<=0;
   42607: out<=1;
   42608: out<=1;
   42609: out<=0;
   42610: out<=0;
   42611: out<=1;
   42612: out<=1;
   42613: out<=1;
   42614: out<=1;
   42615: out<=1;
   42616: out<=1;
   42617: out<=1;
   42618: out<=0;
   42619: out<=0;
   42620: out<=1;
   42621: out<=0;
   42622: out<=1;
   42623: out<=0;
   42624: out<=1;
   42625: out<=0;
   42626: out<=0;
   42627: out<=1;
   42628: out<=1;
   42629: out<=1;
   42630: out<=1;
   42631: out<=1;
   42632: out<=1;
   42633: out<=1;
   42634: out<=0;
   42635: out<=0;
   42636: out<=1;
   42637: out<=0;
   42638: out<=1;
   42639: out<=0;
   42640: out<=0;
   42641: out<=1;
   42642: out<=1;
   42643: out<=0;
   42644: out<=0;
   42645: out<=0;
   42646: out<=0;
   42647: out<=0;
   42648: out<=0;
   42649: out<=0;
   42650: out<=1;
   42651: out<=1;
   42652: out<=0;
   42653: out<=1;
   42654: out<=0;
   42655: out<=1;
   42656: out<=1;
   42657: out<=0;
   42658: out<=0;
   42659: out<=1;
   42660: out<=1;
   42661: out<=1;
   42662: out<=1;
   42663: out<=1;
   42664: out<=1;
   42665: out<=1;
   42666: out<=0;
   42667: out<=0;
   42668: out<=1;
   42669: out<=0;
   42670: out<=1;
   42671: out<=0;
   42672: out<=0;
   42673: out<=1;
   42674: out<=1;
   42675: out<=0;
   42676: out<=0;
   42677: out<=0;
   42678: out<=0;
   42679: out<=0;
   42680: out<=0;
   42681: out<=0;
   42682: out<=1;
   42683: out<=1;
   42684: out<=0;
   42685: out<=1;
   42686: out<=0;
   42687: out<=1;
   42688: out<=1;
   42689: out<=0;
   42690: out<=0;
   42691: out<=1;
   42692: out<=1;
   42693: out<=1;
   42694: out<=1;
   42695: out<=1;
   42696: out<=1;
   42697: out<=1;
   42698: out<=0;
   42699: out<=0;
   42700: out<=1;
   42701: out<=0;
   42702: out<=1;
   42703: out<=0;
   42704: out<=1;
   42705: out<=0;
   42706: out<=0;
   42707: out<=1;
   42708: out<=1;
   42709: out<=1;
   42710: out<=1;
   42711: out<=1;
   42712: out<=1;
   42713: out<=1;
   42714: out<=0;
   42715: out<=0;
   42716: out<=1;
   42717: out<=0;
   42718: out<=1;
   42719: out<=0;
   42720: out<=0;
   42721: out<=1;
   42722: out<=1;
   42723: out<=0;
   42724: out<=0;
   42725: out<=0;
   42726: out<=0;
   42727: out<=0;
   42728: out<=0;
   42729: out<=0;
   42730: out<=1;
   42731: out<=1;
   42732: out<=0;
   42733: out<=1;
   42734: out<=0;
   42735: out<=1;
   42736: out<=0;
   42737: out<=1;
   42738: out<=1;
   42739: out<=0;
   42740: out<=0;
   42741: out<=0;
   42742: out<=0;
   42743: out<=0;
   42744: out<=0;
   42745: out<=0;
   42746: out<=1;
   42747: out<=1;
   42748: out<=0;
   42749: out<=1;
   42750: out<=0;
   42751: out<=1;
   42752: out<=0;
   42753: out<=0;
   42754: out<=0;
   42755: out<=0;
   42756: out<=1;
   42757: out<=0;
   42758: out<=0;
   42759: out<=1;
   42760: out<=1;
   42761: out<=0;
   42762: out<=1;
   42763: out<=0;
   42764: out<=0;
   42765: out<=0;
   42766: out<=1;
   42767: out<=1;
   42768: out<=1;
   42769: out<=1;
   42770: out<=1;
   42771: out<=1;
   42772: out<=0;
   42773: out<=1;
   42774: out<=1;
   42775: out<=0;
   42776: out<=0;
   42777: out<=1;
   42778: out<=0;
   42779: out<=1;
   42780: out<=1;
   42781: out<=1;
   42782: out<=0;
   42783: out<=0;
   42784: out<=1;
   42785: out<=1;
   42786: out<=1;
   42787: out<=1;
   42788: out<=0;
   42789: out<=1;
   42790: out<=1;
   42791: out<=0;
   42792: out<=0;
   42793: out<=1;
   42794: out<=0;
   42795: out<=1;
   42796: out<=1;
   42797: out<=1;
   42798: out<=0;
   42799: out<=0;
   42800: out<=0;
   42801: out<=0;
   42802: out<=0;
   42803: out<=0;
   42804: out<=1;
   42805: out<=0;
   42806: out<=0;
   42807: out<=1;
   42808: out<=1;
   42809: out<=0;
   42810: out<=1;
   42811: out<=0;
   42812: out<=0;
   42813: out<=0;
   42814: out<=1;
   42815: out<=1;
   42816: out<=0;
   42817: out<=0;
   42818: out<=0;
   42819: out<=0;
   42820: out<=1;
   42821: out<=0;
   42822: out<=0;
   42823: out<=1;
   42824: out<=1;
   42825: out<=0;
   42826: out<=1;
   42827: out<=0;
   42828: out<=0;
   42829: out<=0;
   42830: out<=1;
   42831: out<=1;
   42832: out<=0;
   42833: out<=0;
   42834: out<=0;
   42835: out<=0;
   42836: out<=1;
   42837: out<=0;
   42838: out<=0;
   42839: out<=1;
   42840: out<=1;
   42841: out<=0;
   42842: out<=1;
   42843: out<=0;
   42844: out<=0;
   42845: out<=0;
   42846: out<=1;
   42847: out<=1;
   42848: out<=0;
   42849: out<=0;
   42850: out<=0;
   42851: out<=0;
   42852: out<=1;
   42853: out<=0;
   42854: out<=0;
   42855: out<=1;
   42856: out<=1;
   42857: out<=0;
   42858: out<=1;
   42859: out<=0;
   42860: out<=0;
   42861: out<=0;
   42862: out<=1;
   42863: out<=1;
   42864: out<=0;
   42865: out<=0;
   42866: out<=0;
   42867: out<=0;
   42868: out<=1;
   42869: out<=0;
   42870: out<=0;
   42871: out<=1;
   42872: out<=1;
   42873: out<=0;
   42874: out<=1;
   42875: out<=0;
   42876: out<=0;
   42877: out<=0;
   42878: out<=1;
   42879: out<=1;
   42880: out<=0;
   42881: out<=0;
   42882: out<=0;
   42883: out<=0;
   42884: out<=1;
   42885: out<=0;
   42886: out<=0;
   42887: out<=1;
   42888: out<=1;
   42889: out<=0;
   42890: out<=1;
   42891: out<=0;
   42892: out<=0;
   42893: out<=0;
   42894: out<=1;
   42895: out<=1;
   42896: out<=0;
   42897: out<=0;
   42898: out<=0;
   42899: out<=0;
   42900: out<=1;
   42901: out<=0;
   42902: out<=0;
   42903: out<=1;
   42904: out<=1;
   42905: out<=0;
   42906: out<=1;
   42907: out<=0;
   42908: out<=0;
   42909: out<=0;
   42910: out<=1;
   42911: out<=1;
   42912: out<=1;
   42913: out<=1;
   42914: out<=1;
   42915: out<=1;
   42916: out<=0;
   42917: out<=1;
   42918: out<=1;
   42919: out<=0;
   42920: out<=0;
   42921: out<=1;
   42922: out<=0;
   42923: out<=1;
   42924: out<=1;
   42925: out<=1;
   42926: out<=0;
   42927: out<=0;
   42928: out<=1;
   42929: out<=1;
   42930: out<=1;
   42931: out<=1;
   42932: out<=0;
   42933: out<=1;
   42934: out<=1;
   42935: out<=0;
   42936: out<=0;
   42937: out<=1;
   42938: out<=0;
   42939: out<=1;
   42940: out<=1;
   42941: out<=1;
   42942: out<=0;
   42943: out<=0;
   42944: out<=0;
   42945: out<=0;
   42946: out<=0;
   42947: out<=0;
   42948: out<=1;
   42949: out<=0;
   42950: out<=0;
   42951: out<=1;
   42952: out<=1;
   42953: out<=0;
   42954: out<=1;
   42955: out<=0;
   42956: out<=0;
   42957: out<=0;
   42958: out<=1;
   42959: out<=1;
   42960: out<=1;
   42961: out<=1;
   42962: out<=1;
   42963: out<=1;
   42964: out<=0;
   42965: out<=1;
   42966: out<=1;
   42967: out<=0;
   42968: out<=0;
   42969: out<=1;
   42970: out<=0;
   42971: out<=1;
   42972: out<=1;
   42973: out<=1;
   42974: out<=0;
   42975: out<=0;
   42976: out<=0;
   42977: out<=0;
   42978: out<=0;
   42979: out<=0;
   42980: out<=1;
   42981: out<=0;
   42982: out<=0;
   42983: out<=1;
   42984: out<=1;
   42985: out<=0;
   42986: out<=1;
   42987: out<=0;
   42988: out<=0;
   42989: out<=0;
   42990: out<=1;
   42991: out<=1;
   42992: out<=1;
   42993: out<=1;
   42994: out<=1;
   42995: out<=1;
   42996: out<=0;
   42997: out<=1;
   42998: out<=1;
   42999: out<=0;
   43000: out<=0;
   43001: out<=1;
   43002: out<=0;
   43003: out<=1;
   43004: out<=1;
   43005: out<=1;
   43006: out<=0;
   43007: out<=0;
   43008: out<=0;
   43009: out<=0;
   43010: out<=0;
   43011: out<=0;
   43012: out<=1;
   43013: out<=0;
   43014: out<=0;
   43015: out<=1;
   43016: out<=0;
   43017: out<=1;
   43018: out<=0;
   43019: out<=1;
   43020: out<=1;
   43021: out<=1;
   43022: out<=0;
   43023: out<=0;
   43024: out<=1;
   43025: out<=1;
   43026: out<=1;
   43027: out<=1;
   43028: out<=0;
   43029: out<=1;
   43030: out<=1;
   43031: out<=0;
   43032: out<=1;
   43033: out<=0;
   43034: out<=1;
   43035: out<=0;
   43036: out<=0;
   43037: out<=0;
   43038: out<=1;
   43039: out<=1;
   43040: out<=0;
   43041: out<=0;
   43042: out<=0;
   43043: out<=0;
   43044: out<=1;
   43045: out<=0;
   43046: out<=0;
   43047: out<=1;
   43048: out<=0;
   43049: out<=1;
   43050: out<=0;
   43051: out<=1;
   43052: out<=1;
   43053: out<=1;
   43054: out<=0;
   43055: out<=0;
   43056: out<=1;
   43057: out<=1;
   43058: out<=1;
   43059: out<=1;
   43060: out<=0;
   43061: out<=1;
   43062: out<=1;
   43063: out<=0;
   43064: out<=1;
   43065: out<=0;
   43066: out<=1;
   43067: out<=0;
   43068: out<=0;
   43069: out<=0;
   43070: out<=1;
   43071: out<=1;
   43072: out<=0;
   43073: out<=0;
   43074: out<=0;
   43075: out<=0;
   43076: out<=1;
   43077: out<=0;
   43078: out<=0;
   43079: out<=1;
   43080: out<=0;
   43081: out<=1;
   43082: out<=0;
   43083: out<=1;
   43084: out<=1;
   43085: out<=1;
   43086: out<=0;
   43087: out<=0;
   43088: out<=0;
   43089: out<=0;
   43090: out<=0;
   43091: out<=0;
   43092: out<=1;
   43093: out<=0;
   43094: out<=0;
   43095: out<=1;
   43096: out<=0;
   43097: out<=1;
   43098: out<=0;
   43099: out<=1;
   43100: out<=1;
   43101: out<=1;
   43102: out<=0;
   43103: out<=0;
   43104: out<=1;
   43105: out<=1;
   43106: out<=1;
   43107: out<=1;
   43108: out<=0;
   43109: out<=1;
   43110: out<=1;
   43111: out<=0;
   43112: out<=1;
   43113: out<=0;
   43114: out<=1;
   43115: out<=0;
   43116: out<=0;
   43117: out<=0;
   43118: out<=1;
   43119: out<=1;
   43120: out<=1;
   43121: out<=1;
   43122: out<=1;
   43123: out<=1;
   43124: out<=0;
   43125: out<=1;
   43126: out<=1;
   43127: out<=0;
   43128: out<=1;
   43129: out<=0;
   43130: out<=1;
   43131: out<=0;
   43132: out<=0;
   43133: out<=0;
   43134: out<=1;
   43135: out<=1;
   43136: out<=0;
   43137: out<=0;
   43138: out<=0;
   43139: out<=0;
   43140: out<=1;
   43141: out<=0;
   43142: out<=0;
   43143: out<=1;
   43144: out<=0;
   43145: out<=1;
   43146: out<=0;
   43147: out<=1;
   43148: out<=1;
   43149: out<=1;
   43150: out<=0;
   43151: out<=0;
   43152: out<=0;
   43153: out<=0;
   43154: out<=0;
   43155: out<=0;
   43156: out<=1;
   43157: out<=0;
   43158: out<=0;
   43159: out<=1;
   43160: out<=0;
   43161: out<=1;
   43162: out<=0;
   43163: out<=1;
   43164: out<=1;
   43165: out<=1;
   43166: out<=0;
   43167: out<=0;
   43168: out<=0;
   43169: out<=0;
   43170: out<=0;
   43171: out<=0;
   43172: out<=1;
   43173: out<=0;
   43174: out<=0;
   43175: out<=1;
   43176: out<=0;
   43177: out<=1;
   43178: out<=0;
   43179: out<=1;
   43180: out<=1;
   43181: out<=1;
   43182: out<=0;
   43183: out<=0;
   43184: out<=0;
   43185: out<=0;
   43186: out<=0;
   43187: out<=0;
   43188: out<=1;
   43189: out<=0;
   43190: out<=0;
   43191: out<=1;
   43192: out<=0;
   43193: out<=1;
   43194: out<=0;
   43195: out<=1;
   43196: out<=1;
   43197: out<=1;
   43198: out<=0;
   43199: out<=0;
   43200: out<=0;
   43201: out<=0;
   43202: out<=0;
   43203: out<=0;
   43204: out<=1;
   43205: out<=0;
   43206: out<=0;
   43207: out<=1;
   43208: out<=0;
   43209: out<=1;
   43210: out<=0;
   43211: out<=1;
   43212: out<=1;
   43213: out<=1;
   43214: out<=0;
   43215: out<=0;
   43216: out<=1;
   43217: out<=1;
   43218: out<=1;
   43219: out<=1;
   43220: out<=0;
   43221: out<=1;
   43222: out<=1;
   43223: out<=0;
   43224: out<=1;
   43225: out<=0;
   43226: out<=1;
   43227: out<=0;
   43228: out<=0;
   43229: out<=0;
   43230: out<=1;
   43231: out<=1;
   43232: out<=1;
   43233: out<=1;
   43234: out<=1;
   43235: out<=1;
   43236: out<=0;
   43237: out<=1;
   43238: out<=1;
   43239: out<=0;
   43240: out<=1;
   43241: out<=0;
   43242: out<=1;
   43243: out<=0;
   43244: out<=0;
   43245: out<=0;
   43246: out<=1;
   43247: out<=1;
   43248: out<=0;
   43249: out<=0;
   43250: out<=0;
   43251: out<=0;
   43252: out<=1;
   43253: out<=0;
   43254: out<=0;
   43255: out<=1;
   43256: out<=0;
   43257: out<=1;
   43258: out<=0;
   43259: out<=1;
   43260: out<=1;
   43261: out<=1;
   43262: out<=0;
   43263: out<=0;
   43264: out<=1;
   43265: out<=0;
   43266: out<=0;
   43267: out<=1;
   43268: out<=1;
   43269: out<=1;
   43270: out<=1;
   43271: out<=1;
   43272: out<=0;
   43273: out<=0;
   43274: out<=1;
   43275: out<=1;
   43276: out<=0;
   43277: out<=1;
   43278: out<=0;
   43279: out<=1;
   43280: out<=1;
   43281: out<=0;
   43282: out<=0;
   43283: out<=1;
   43284: out<=1;
   43285: out<=1;
   43286: out<=1;
   43287: out<=1;
   43288: out<=0;
   43289: out<=0;
   43290: out<=1;
   43291: out<=1;
   43292: out<=0;
   43293: out<=1;
   43294: out<=0;
   43295: out<=1;
   43296: out<=0;
   43297: out<=1;
   43298: out<=1;
   43299: out<=0;
   43300: out<=0;
   43301: out<=0;
   43302: out<=0;
   43303: out<=0;
   43304: out<=1;
   43305: out<=1;
   43306: out<=0;
   43307: out<=0;
   43308: out<=1;
   43309: out<=0;
   43310: out<=1;
   43311: out<=0;
   43312: out<=0;
   43313: out<=1;
   43314: out<=1;
   43315: out<=0;
   43316: out<=0;
   43317: out<=0;
   43318: out<=0;
   43319: out<=0;
   43320: out<=1;
   43321: out<=1;
   43322: out<=0;
   43323: out<=0;
   43324: out<=1;
   43325: out<=0;
   43326: out<=1;
   43327: out<=0;
   43328: out<=1;
   43329: out<=0;
   43330: out<=0;
   43331: out<=1;
   43332: out<=1;
   43333: out<=1;
   43334: out<=1;
   43335: out<=1;
   43336: out<=0;
   43337: out<=0;
   43338: out<=1;
   43339: out<=1;
   43340: out<=0;
   43341: out<=1;
   43342: out<=0;
   43343: out<=1;
   43344: out<=0;
   43345: out<=1;
   43346: out<=1;
   43347: out<=0;
   43348: out<=0;
   43349: out<=0;
   43350: out<=0;
   43351: out<=0;
   43352: out<=1;
   43353: out<=1;
   43354: out<=0;
   43355: out<=0;
   43356: out<=1;
   43357: out<=0;
   43358: out<=1;
   43359: out<=0;
   43360: out<=1;
   43361: out<=0;
   43362: out<=0;
   43363: out<=1;
   43364: out<=1;
   43365: out<=1;
   43366: out<=1;
   43367: out<=1;
   43368: out<=0;
   43369: out<=0;
   43370: out<=1;
   43371: out<=1;
   43372: out<=0;
   43373: out<=1;
   43374: out<=0;
   43375: out<=1;
   43376: out<=0;
   43377: out<=1;
   43378: out<=1;
   43379: out<=0;
   43380: out<=0;
   43381: out<=0;
   43382: out<=0;
   43383: out<=0;
   43384: out<=1;
   43385: out<=1;
   43386: out<=0;
   43387: out<=0;
   43388: out<=1;
   43389: out<=0;
   43390: out<=1;
   43391: out<=0;
   43392: out<=1;
   43393: out<=0;
   43394: out<=0;
   43395: out<=1;
   43396: out<=1;
   43397: out<=1;
   43398: out<=1;
   43399: out<=1;
   43400: out<=0;
   43401: out<=0;
   43402: out<=1;
   43403: out<=1;
   43404: out<=0;
   43405: out<=1;
   43406: out<=0;
   43407: out<=1;
   43408: out<=0;
   43409: out<=1;
   43410: out<=1;
   43411: out<=0;
   43412: out<=0;
   43413: out<=0;
   43414: out<=0;
   43415: out<=0;
   43416: out<=1;
   43417: out<=1;
   43418: out<=0;
   43419: out<=0;
   43420: out<=1;
   43421: out<=0;
   43422: out<=1;
   43423: out<=0;
   43424: out<=0;
   43425: out<=1;
   43426: out<=1;
   43427: out<=0;
   43428: out<=0;
   43429: out<=0;
   43430: out<=0;
   43431: out<=0;
   43432: out<=1;
   43433: out<=1;
   43434: out<=0;
   43435: out<=0;
   43436: out<=1;
   43437: out<=0;
   43438: out<=1;
   43439: out<=0;
   43440: out<=1;
   43441: out<=0;
   43442: out<=0;
   43443: out<=1;
   43444: out<=1;
   43445: out<=1;
   43446: out<=1;
   43447: out<=1;
   43448: out<=0;
   43449: out<=0;
   43450: out<=1;
   43451: out<=1;
   43452: out<=0;
   43453: out<=1;
   43454: out<=0;
   43455: out<=1;
   43456: out<=1;
   43457: out<=0;
   43458: out<=0;
   43459: out<=1;
   43460: out<=1;
   43461: out<=1;
   43462: out<=1;
   43463: out<=1;
   43464: out<=0;
   43465: out<=0;
   43466: out<=1;
   43467: out<=1;
   43468: out<=0;
   43469: out<=1;
   43470: out<=0;
   43471: out<=1;
   43472: out<=1;
   43473: out<=0;
   43474: out<=0;
   43475: out<=1;
   43476: out<=1;
   43477: out<=1;
   43478: out<=1;
   43479: out<=1;
   43480: out<=0;
   43481: out<=0;
   43482: out<=1;
   43483: out<=1;
   43484: out<=0;
   43485: out<=1;
   43486: out<=0;
   43487: out<=1;
   43488: out<=1;
   43489: out<=0;
   43490: out<=0;
   43491: out<=1;
   43492: out<=1;
   43493: out<=1;
   43494: out<=1;
   43495: out<=1;
   43496: out<=0;
   43497: out<=0;
   43498: out<=1;
   43499: out<=1;
   43500: out<=0;
   43501: out<=1;
   43502: out<=0;
   43503: out<=1;
   43504: out<=1;
   43505: out<=0;
   43506: out<=0;
   43507: out<=1;
   43508: out<=1;
   43509: out<=1;
   43510: out<=1;
   43511: out<=1;
   43512: out<=0;
   43513: out<=0;
   43514: out<=1;
   43515: out<=1;
   43516: out<=0;
   43517: out<=1;
   43518: out<=0;
   43519: out<=1;
   43520: out<=0;
   43521: out<=1;
   43522: out<=0;
   43523: out<=1;
   43524: out<=0;
   43525: out<=0;
   43526: out<=1;
   43527: out<=1;
   43528: out<=0;
   43529: out<=0;
   43530: out<=0;
   43531: out<=0;
   43532: out<=0;
   43533: out<=1;
   43534: out<=1;
   43535: out<=0;
   43536: out<=0;
   43537: out<=1;
   43538: out<=0;
   43539: out<=1;
   43540: out<=0;
   43541: out<=0;
   43542: out<=1;
   43543: out<=1;
   43544: out<=0;
   43545: out<=0;
   43546: out<=0;
   43547: out<=0;
   43548: out<=0;
   43549: out<=1;
   43550: out<=1;
   43551: out<=0;
   43552: out<=0;
   43553: out<=1;
   43554: out<=0;
   43555: out<=1;
   43556: out<=0;
   43557: out<=0;
   43558: out<=1;
   43559: out<=1;
   43560: out<=0;
   43561: out<=0;
   43562: out<=0;
   43563: out<=0;
   43564: out<=0;
   43565: out<=1;
   43566: out<=1;
   43567: out<=0;
   43568: out<=0;
   43569: out<=1;
   43570: out<=0;
   43571: out<=1;
   43572: out<=0;
   43573: out<=0;
   43574: out<=1;
   43575: out<=1;
   43576: out<=0;
   43577: out<=0;
   43578: out<=0;
   43579: out<=0;
   43580: out<=0;
   43581: out<=1;
   43582: out<=1;
   43583: out<=0;
   43584: out<=0;
   43585: out<=1;
   43586: out<=0;
   43587: out<=1;
   43588: out<=0;
   43589: out<=0;
   43590: out<=1;
   43591: out<=1;
   43592: out<=0;
   43593: out<=0;
   43594: out<=0;
   43595: out<=0;
   43596: out<=0;
   43597: out<=1;
   43598: out<=1;
   43599: out<=0;
   43600: out<=1;
   43601: out<=0;
   43602: out<=1;
   43603: out<=0;
   43604: out<=1;
   43605: out<=1;
   43606: out<=0;
   43607: out<=0;
   43608: out<=1;
   43609: out<=1;
   43610: out<=1;
   43611: out<=1;
   43612: out<=1;
   43613: out<=0;
   43614: out<=0;
   43615: out<=1;
   43616: out<=1;
   43617: out<=0;
   43618: out<=1;
   43619: out<=0;
   43620: out<=1;
   43621: out<=1;
   43622: out<=0;
   43623: out<=0;
   43624: out<=1;
   43625: out<=1;
   43626: out<=1;
   43627: out<=1;
   43628: out<=1;
   43629: out<=0;
   43630: out<=0;
   43631: out<=1;
   43632: out<=0;
   43633: out<=1;
   43634: out<=0;
   43635: out<=1;
   43636: out<=0;
   43637: out<=0;
   43638: out<=1;
   43639: out<=1;
   43640: out<=0;
   43641: out<=0;
   43642: out<=0;
   43643: out<=0;
   43644: out<=0;
   43645: out<=1;
   43646: out<=1;
   43647: out<=0;
   43648: out<=0;
   43649: out<=1;
   43650: out<=0;
   43651: out<=1;
   43652: out<=0;
   43653: out<=0;
   43654: out<=1;
   43655: out<=1;
   43656: out<=0;
   43657: out<=0;
   43658: out<=0;
   43659: out<=0;
   43660: out<=0;
   43661: out<=1;
   43662: out<=1;
   43663: out<=0;
   43664: out<=1;
   43665: out<=0;
   43666: out<=1;
   43667: out<=0;
   43668: out<=1;
   43669: out<=1;
   43670: out<=0;
   43671: out<=0;
   43672: out<=1;
   43673: out<=1;
   43674: out<=1;
   43675: out<=1;
   43676: out<=1;
   43677: out<=0;
   43678: out<=0;
   43679: out<=1;
   43680: out<=0;
   43681: out<=1;
   43682: out<=0;
   43683: out<=1;
   43684: out<=0;
   43685: out<=0;
   43686: out<=1;
   43687: out<=1;
   43688: out<=0;
   43689: out<=0;
   43690: out<=0;
   43691: out<=0;
   43692: out<=0;
   43693: out<=1;
   43694: out<=1;
   43695: out<=0;
   43696: out<=1;
   43697: out<=0;
   43698: out<=1;
   43699: out<=0;
   43700: out<=1;
   43701: out<=1;
   43702: out<=0;
   43703: out<=0;
   43704: out<=1;
   43705: out<=1;
   43706: out<=1;
   43707: out<=1;
   43708: out<=1;
   43709: out<=0;
   43710: out<=0;
   43711: out<=1;
   43712: out<=0;
   43713: out<=1;
   43714: out<=0;
   43715: out<=1;
   43716: out<=0;
   43717: out<=0;
   43718: out<=1;
   43719: out<=1;
   43720: out<=0;
   43721: out<=0;
   43722: out<=0;
   43723: out<=0;
   43724: out<=0;
   43725: out<=1;
   43726: out<=1;
   43727: out<=0;
   43728: out<=0;
   43729: out<=1;
   43730: out<=0;
   43731: out<=1;
   43732: out<=0;
   43733: out<=0;
   43734: out<=1;
   43735: out<=1;
   43736: out<=0;
   43737: out<=0;
   43738: out<=0;
   43739: out<=0;
   43740: out<=0;
   43741: out<=1;
   43742: out<=1;
   43743: out<=0;
   43744: out<=1;
   43745: out<=0;
   43746: out<=1;
   43747: out<=0;
   43748: out<=1;
   43749: out<=1;
   43750: out<=0;
   43751: out<=0;
   43752: out<=1;
   43753: out<=1;
   43754: out<=1;
   43755: out<=1;
   43756: out<=1;
   43757: out<=0;
   43758: out<=0;
   43759: out<=1;
   43760: out<=1;
   43761: out<=0;
   43762: out<=1;
   43763: out<=0;
   43764: out<=1;
   43765: out<=1;
   43766: out<=0;
   43767: out<=0;
   43768: out<=1;
   43769: out<=1;
   43770: out<=1;
   43771: out<=1;
   43772: out<=1;
   43773: out<=0;
   43774: out<=0;
   43775: out<=1;
   43776: out<=1;
   43777: out<=1;
   43778: out<=0;
   43779: out<=0;
   43780: out<=0;
   43781: out<=1;
   43782: out<=0;
   43783: out<=1;
   43784: out<=0;
   43785: out<=1;
   43786: out<=1;
   43787: out<=0;
   43788: out<=1;
   43789: out<=1;
   43790: out<=1;
   43791: out<=1;
   43792: out<=0;
   43793: out<=0;
   43794: out<=1;
   43795: out<=1;
   43796: out<=1;
   43797: out<=0;
   43798: out<=1;
   43799: out<=0;
   43800: out<=1;
   43801: out<=0;
   43802: out<=0;
   43803: out<=1;
   43804: out<=0;
   43805: out<=0;
   43806: out<=0;
   43807: out<=0;
   43808: out<=0;
   43809: out<=0;
   43810: out<=1;
   43811: out<=1;
   43812: out<=1;
   43813: out<=0;
   43814: out<=1;
   43815: out<=0;
   43816: out<=1;
   43817: out<=0;
   43818: out<=0;
   43819: out<=1;
   43820: out<=0;
   43821: out<=0;
   43822: out<=0;
   43823: out<=0;
   43824: out<=1;
   43825: out<=1;
   43826: out<=0;
   43827: out<=0;
   43828: out<=0;
   43829: out<=1;
   43830: out<=0;
   43831: out<=1;
   43832: out<=0;
   43833: out<=1;
   43834: out<=1;
   43835: out<=0;
   43836: out<=1;
   43837: out<=1;
   43838: out<=1;
   43839: out<=1;
   43840: out<=1;
   43841: out<=1;
   43842: out<=0;
   43843: out<=0;
   43844: out<=0;
   43845: out<=1;
   43846: out<=0;
   43847: out<=1;
   43848: out<=0;
   43849: out<=1;
   43850: out<=1;
   43851: out<=0;
   43852: out<=1;
   43853: out<=1;
   43854: out<=1;
   43855: out<=1;
   43856: out<=1;
   43857: out<=1;
   43858: out<=0;
   43859: out<=0;
   43860: out<=0;
   43861: out<=1;
   43862: out<=0;
   43863: out<=1;
   43864: out<=0;
   43865: out<=1;
   43866: out<=1;
   43867: out<=0;
   43868: out<=1;
   43869: out<=1;
   43870: out<=1;
   43871: out<=1;
   43872: out<=1;
   43873: out<=1;
   43874: out<=0;
   43875: out<=0;
   43876: out<=0;
   43877: out<=1;
   43878: out<=0;
   43879: out<=1;
   43880: out<=0;
   43881: out<=1;
   43882: out<=1;
   43883: out<=0;
   43884: out<=1;
   43885: out<=1;
   43886: out<=1;
   43887: out<=1;
   43888: out<=1;
   43889: out<=1;
   43890: out<=0;
   43891: out<=0;
   43892: out<=0;
   43893: out<=1;
   43894: out<=0;
   43895: out<=1;
   43896: out<=0;
   43897: out<=1;
   43898: out<=1;
   43899: out<=0;
   43900: out<=1;
   43901: out<=1;
   43902: out<=1;
   43903: out<=1;
   43904: out<=1;
   43905: out<=1;
   43906: out<=0;
   43907: out<=0;
   43908: out<=0;
   43909: out<=1;
   43910: out<=0;
   43911: out<=1;
   43912: out<=0;
   43913: out<=1;
   43914: out<=1;
   43915: out<=0;
   43916: out<=1;
   43917: out<=1;
   43918: out<=1;
   43919: out<=1;
   43920: out<=1;
   43921: out<=1;
   43922: out<=0;
   43923: out<=0;
   43924: out<=0;
   43925: out<=1;
   43926: out<=0;
   43927: out<=1;
   43928: out<=0;
   43929: out<=1;
   43930: out<=1;
   43931: out<=0;
   43932: out<=1;
   43933: out<=1;
   43934: out<=1;
   43935: out<=1;
   43936: out<=0;
   43937: out<=0;
   43938: out<=1;
   43939: out<=1;
   43940: out<=1;
   43941: out<=0;
   43942: out<=1;
   43943: out<=0;
   43944: out<=1;
   43945: out<=0;
   43946: out<=0;
   43947: out<=1;
   43948: out<=0;
   43949: out<=0;
   43950: out<=0;
   43951: out<=0;
   43952: out<=0;
   43953: out<=0;
   43954: out<=1;
   43955: out<=1;
   43956: out<=1;
   43957: out<=0;
   43958: out<=1;
   43959: out<=0;
   43960: out<=1;
   43961: out<=0;
   43962: out<=0;
   43963: out<=1;
   43964: out<=0;
   43965: out<=0;
   43966: out<=0;
   43967: out<=0;
   43968: out<=1;
   43969: out<=1;
   43970: out<=0;
   43971: out<=0;
   43972: out<=0;
   43973: out<=1;
   43974: out<=0;
   43975: out<=1;
   43976: out<=0;
   43977: out<=1;
   43978: out<=1;
   43979: out<=0;
   43980: out<=1;
   43981: out<=1;
   43982: out<=1;
   43983: out<=1;
   43984: out<=0;
   43985: out<=0;
   43986: out<=1;
   43987: out<=1;
   43988: out<=1;
   43989: out<=0;
   43990: out<=1;
   43991: out<=0;
   43992: out<=1;
   43993: out<=0;
   43994: out<=0;
   43995: out<=1;
   43996: out<=0;
   43997: out<=0;
   43998: out<=0;
   43999: out<=0;
   44000: out<=1;
   44001: out<=1;
   44002: out<=0;
   44003: out<=0;
   44004: out<=0;
   44005: out<=1;
   44006: out<=0;
   44007: out<=1;
   44008: out<=0;
   44009: out<=1;
   44010: out<=1;
   44011: out<=0;
   44012: out<=1;
   44013: out<=1;
   44014: out<=1;
   44015: out<=1;
   44016: out<=0;
   44017: out<=0;
   44018: out<=1;
   44019: out<=1;
   44020: out<=1;
   44021: out<=0;
   44022: out<=1;
   44023: out<=0;
   44024: out<=1;
   44025: out<=0;
   44026: out<=0;
   44027: out<=1;
   44028: out<=0;
   44029: out<=0;
   44030: out<=0;
   44031: out<=0;
   44032: out<=0;
   44033: out<=1;
   44034: out<=1;
   44035: out<=0;
   44036: out<=1;
   44037: out<=1;
   44038: out<=1;
   44039: out<=1;
   44040: out<=0;
   44041: out<=0;
   44042: out<=1;
   44043: out<=1;
   44044: out<=1;
   44045: out<=0;
   44046: out<=1;
   44047: out<=0;
   44048: out<=1;
   44049: out<=0;
   44050: out<=0;
   44051: out<=1;
   44052: out<=0;
   44053: out<=0;
   44054: out<=0;
   44055: out<=0;
   44056: out<=1;
   44057: out<=1;
   44058: out<=0;
   44059: out<=0;
   44060: out<=0;
   44061: out<=1;
   44062: out<=0;
   44063: out<=1;
   44064: out<=0;
   44065: out<=1;
   44066: out<=1;
   44067: out<=0;
   44068: out<=1;
   44069: out<=1;
   44070: out<=1;
   44071: out<=1;
   44072: out<=0;
   44073: out<=0;
   44074: out<=1;
   44075: out<=1;
   44076: out<=1;
   44077: out<=0;
   44078: out<=1;
   44079: out<=0;
   44080: out<=1;
   44081: out<=0;
   44082: out<=0;
   44083: out<=1;
   44084: out<=0;
   44085: out<=0;
   44086: out<=0;
   44087: out<=0;
   44088: out<=1;
   44089: out<=1;
   44090: out<=0;
   44091: out<=0;
   44092: out<=0;
   44093: out<=1;
   44094: out<=0;
   44095: out<=1;
   44096: out<=0;
   44097: out<=1;
   44098: out<=1;
   44099: out<=0;
   44100: out<=1;
   44101: out<=1;
   44102: out<=1;
   44103: out<=1;
   44104: out<=0;
   44105: out<=0;
   44106: out<=1;
   44107: out<=1;
   44108: out<=1;
   44109: out<=0;
   44110: out<=1;
   44111: out<=0;
   44112: out<=0;
   44113: out<=1;
   44114: out<=1;
   44115: out<=0;
   44116: out<=1;
   44117: out<=1;
   44118: out<=1;
   44119: out<=1;
   44120: out<=0;
   44121: out<=0;
   44122: out<=1;
   44123: out<=1;
   44124: out<=1;
   44125: out<=0;
   44126: out<=1;
   44127: out<=0;
   44128: out<=1;
   44129: out<=0;
   44130: out<=0;
   44131: out<=1;
   44132: out<=0;
   44133: out<=0;
   44134: out<=0;
   44135: out<=0;
   44136: out<=1;
   44137: out<=1;
   44138: out<=0;
   44139: out<=0;
   44140: out<=0;
   44141: out<=1;
   44142: out<=0;
   44143: out<=1;
   44144: out<=1;
   44145: out<=0;
   44146: out<=0;
   44147: out<=1;
   44148: out<=0;
   44149: out<=0;
   44150: out<=0;
   44151: out<=0;
   44152: out<=1;
   44153: out<=1;
   44154: out<=0;
   44155: out<=0;
   44156: out<=0;
   44157: out<=1;
   44158: out<=0;
   44159: out<=1;
   44160: out<=0;
   44161: out<=1;
   44162: out<=1;
   44163: out<=0;
   44164: out<=1;
   44165: out<=1;
   44166: out<=1;
   44167: out<=1;
   44168: out<=0;
   44169: out<=0;
   44170: out<=1;
   44171: out<=1;
   44172: out<=1;
   44173: out<=0;
   44174: out<=1;
   44175: out<=0;
   44176: out<=0;
   44177: out<=1;
   44178: out<=1;
   44179: out<=0;
   44180: out<=1;
   44181: out<=1;
   44182: out<=1;
   44183: out<=1;
   44184: out<=0;
   44185: out<=0;
   44186: out<=1;
   44187: out<=1;
   44188: out<=1;
   44189: out<=0;
   44190: out<=1;
   44191: out<=0;
   44192: out<=0;
   44193: out<=1;
   44194: out<=1;
   44195: out<=0;
   44196: out<=1;
   44197: out<=1;
   44198: out<=1;
   44199: out<=1;
   44200: out<=0;
   44201: out<=0;
   44202: out<=1;
   44203: out<=1;
   44204: out<=1;
   44205: out<=0;
   44206: out<=1;
   44207: out<=0;
   44208: out<=0;
   44209: out<=1;
   44210: out<=1;
   44211: out<=0;
   44212: out<=1;
   44213: out<=1;
   44214: out<=1;
   44215: out<=1;
   44216: out<=0;
   44217: out<=0;
   44218: out<=1;
   44219: out<=1;
   44220: out<=1;
   44221: out<=0;
   44222: out<=1;
   44223: out<=0;
   44224: out<=0;
   44225: out<=1;
   44226: out<=1;
   44227: out<=0;
   44228: out<=1;
   44229: out<=1;
   44230: out<=1;
   44231: out<=1;
   44232: out<=0;
   44233: out<=0;
   44234: out<=1;
   44235: out<=1;
   44236: out<=1;
   44237: out<=0;
   44238: out<=1;
   44239: out<=0;
   44240: out<=1;
   44241: out<=0;
   44242: out<=0;
   44243: out<=1;
   44244: out<=0;
   44245: out<=0;
   44246: out<=0;
   44247: out<=0;
   44248: out<=1;
   44249: out<=1;
   44250: out<=0;
   44251: out<=0;
   44252: out<=0;
   44253: out<=1;
   44254: out<=0;
   44255: out<=1;
   44256: out<=1;
   44257: out<=0;
   44258: out<=0;
   44259: out<=1;
   44260: out<=0;
   44261: out<=0;
   44262: out<=0;
   44263: out<=0;
   44264: out<=1;
   44265: out<=1;
   44266: out<=0;
   44267: out<=0;
   44268: out<=0;
   44269: out<=1;
   44270: out<=0;
   44271: out<=1;
   44272: out<=0;
   44273: out<=1;
   44274: out<=1;
   44275: out<=0;
   44276: out<=1;
   44277: out<=1;
   44278: out<=1;
   44279: out<=1;
   44280: out<=0;
   44281: out<=0;
   44282: out<=1;
   44283: out<=1;
   44284: out<=1;
   44285: out<=0;
   44286: out<=1;
   44287: out<=0;
   44288: out<=0;
   44289: out<=0;
   44290: out<=0;
   44291: out<=0;
   44292: out<=0;
   44293: out<=1;
   44294: out<=1;
   44295: out<=0;
   44296: out<=1;
   44297: out<=0;
   44298: out<=1;
   44299: out<=0;
   44300: out<=1;
   44301: out<=1;
   44302: out<=0;
   44303: out<=0;
   44304: out<=0;
   44305: out<=0;
   44306: out<=0;
   44307: out<=0;
   44308: out<=0;
   44309: out<=1;
   44310: out<=1;
   44311: out<=0;
   44312: out<=1;
   44313: out<=0;
   44314: out<=1;
   44315: out<=0;
   44316: out<=1;
   44317: out<=1;
   44318: out<=0;
   44319: out<=0;
   44320: out<=1;
   44321: out<=1;
   44322: out<=1;
   44323: out<=1;
   44324: out<=1;
   44325: out<=0;
   44326: out<=0;
   44327: out<=1;
   44328: out<=0;
   44329: out<=1;
   44330: out<=0;
   44331: out<=1;
   44332: out<=0;
   44333: out<=0;
   44334: out<=1;
   44335: out<=1;
   44336: out<=1;
   44337: out<=1;
   44338: out<=1;
   44339: out<=1;
   44340: out<=1;
   44341: out<=0;
   44342: out<=0;
   44343: out<=1;
   44344: out<=0;
   44345: out<=1;
   44346: out<=0;
   44347: out<=1;
   44348: out<=0;
   44349: out<=0;
   44350: out<=1;
   44351: out<=1;
   44352: out<=0;
   44353: out<=0;
   44354: out<=0;
   44355: out<=0;
   44356: out<=0;
   44357: out<=1;
   44358: out<=1;
   44359: out<=0;
   44360: out<=1;
   44361: out<=0;
   44362: out<=1;
   44363: out<=0;
   44364: out<=1;
   44365: out<=1;
   44366: out<=0;
   44367: out<=0;
   44368: out<=1;
   44369: out<=1;
   44370: out<=1;
   44371: out<=1;
   44372: out<=1;
   44373: out<=0;
   44374: out<=0;
   44375: out<=1;
   44376: out<=0;
   44377: out<=1;
   44378: out<=0;
   44379: out<=1;
   44380: out<=0;
   44381: out<=0;
   44382: out<=1;
   44383: out<=1;
   44384: out<=0;
   44385: out<=0;
   44386: out<=0;
   44387: out<=0;
   44388: out<=0;
   44389: out<=1;
   44390: out<=1;
   44391: out<=0;
   44392: out<=1;
   44393: out<=0;
   44394: out<=1;
   44395: out<=0;
   44396: out<=1;
   44397: out<=1;
   44398: out<=0;
   44399: out<=0;
   44400: out<=1;
   44401: out<=1;
   44402: out<=1;
   44403: out<=1;
   44404: out<=1;
   44405: out<=0;
   44406: out<=0;
   44407: out<=1;
   44408: out<=0;
   44409: out<=1;
   44410: out<=0;
   44411: out<=1;
   44412: out<=0;
   44413: out<=0;
   44414: out<=1;
   44415: out<=1;
   44416: out<=0;
   44417: out<=0;
   44418: out<=0;
   44419: out<=0;
   44420: out<=0;
   44421: out<=1;
   44422: out<=1;
   44423: out<=0;
   44424: out<=1;
   44425: out<=0;
   44426: out<=1;
   44427: out<=0;
   44428: out<=1;
   44429: out<=1;
   44430: out<=0;
   44431: out<=0;
   44432: out<=1;
   44433: out<=1;
   44434: out<=1;
   44435: out<=1;
   44436: out<=1;
   44437: out<=0;
   44438: out<=0;
   44439: out<=1;
   44440: out<=0;
   44441: out<=1;
   44442: out<=0;
   44443: out<=1;
   44444: out<=0;
   44445: out<=0;
   44446: out<=1;
   44447: out<=1;
   44448: out<=1;
   44449: out<=1;
   44450: out<=1;
   44451: out<=1;
   44452: out<=1;
   44453: out<=0;
   44454: out<=0;
   44455: out<=1;
   44456: out<=0;
   44457: out<=1;
   44458: out<=0;
   44459: out<=1;
   44460: out<=0;
   44461: out<=0;
   44462: out<=1;
   44463: out<=1;
   44464: out<=0;
   44465: out<=0;
   44466: out<=0;
   44467: out<=0;
   44468: out<=0;
   44469: out<=1;
   44470: out<=1;
   44471: out<=0;
   44472: out<=1;
   44473: out<=0;
   44474: out<=1;
   44475: out<=0;
   44476: out<=1;
   44477: out<=1;
   44478: out<=0;
   44479: out<=0;
   44480: out<=0;
   44481: out<=0;
   44482: out<=0;
   44483: out<=0;
   44484: out<=0;
   44485: out<=1;
   44486: out<=1;
   44487: out<=0;
   44488: out<=1;
   44489: out<=0;
   44490: out<=1;
   44491: out<=0;
   44492: out<=1;
   44493: out<=1;
   44494: out<=0;
   44495: out<=0;
   44496: out<=0;
   44497: out<=0;
   44498: out<=0;
   44499: out<=0;
   44500: out<=0;
   44501: out<=1;
   44502: out<=1;
   44503: out<=0;
   44504: out<=1;
   44505: out<=0;
   44506: out<=1;
   44507: out<=0;
   44508: out<=1;
   44509: out<=1;
   44510: out<=0;
   44511: out<=0;
   44512: out<=0;
   44513: out<=0;
   44514: out<=0;
   44515: out<=0;
   44516: out<=0;
   44517: out<=1;
   44518: out<=1;
   44519: out<=0;
   44520: out<=1;
   44521: out<=0;
   44522: out<=1;
   44523: out<=0;
   44524: out<=1;
   44525: out<=1;
   44526: out<=0;
   44527: out<=0;
   44528: out<=0;
   44529: out<=0;
   44530: out<=0;
   44531: out<=0;
   44532: out<=0;
   44533: out<=1;
   44534: out<=1;
   44535: out<=0;
   44536: out<=1;
   44537: out<=0;
   44538: out<=1;
   44539: out<=0;
   44540: out<=1;
   44541: out<=1;
   44542: out<=0;
   44543: out<=0;
   44544: out<=1;
   44545: out<=1;
   44546: out<=0;
   44547: out<=0;
   44548: out<=1;
   44549: out<=0;
   44550: out<=1;
   44551: out<=0;
   44552: out<=1;
   44553: out<=0;
   44554: out<=0;
   44555: out<=1;
   44556: out<=1;
   44557: out<=1;
   44558: out<=1;
   44559: out<=1;
   44560: out<=1;
   44561: out<=1;
   44562: out<=0;
   44563: out<=0;
   44564: out<=1;
   44565: out<=0;
   44566: out<=1;
   44567: out<=0;
   44568: out<=1;
   44569: out<=0;
   44570: out<=0;
   44571: out<=1;
   44572: out<=1;
   44573: out<=1;
   44574: out<=1;
   44575: out<=1;
   44576: out<=1;
   44577: out<=1;
   44578: out<=0;
   44579: out<=0;
   44580: out<=1;
   44581: out<=0;
   44582: out<=1;
   44583: out<=0;
   44584: out<=1;
   44585: out<=0;
   44586: out<=0;
   44587: out<=1;
   44588: out<=1;
   44589: out<=1;
   44590: out<=1;
   44591: out<=1;
   44592: out<=1;
   44593: out<=1;
   44594: out<=0;
   44595: out<=0;
   44596: out<=1;
   44597: out<=0;
   44598: out<=1;
   44599: out<=0;
   44600: out<=1;
   44601: out<=0;
   44602: out<=0;
   44603: out<=1;
   44604: out<=1;
   44605: out<=1;
   44606: out<=1;
   44607: out<=1;
   44608: out<=1;
   44609: out<=1;
   44610: out<=0;
   44611: out<=0;
   44612: out<=1;
   44613: out<=0;
   44614: out<=1;
   44615: out<=0;
   44616: out<=1;
   44617: out<=0;
   44618: out<=0;
   44619: out<=1;
   44620: out<=1;
   44621: out<=1;
   44622: out<=1;
   44623: out<=1;
   44624: out<=0;
   44625: out<=0;
   44626: out<=1;
   44627: out<=1;
   44628: out<=0;
   44629: out<=1;
   44630: out<=0;
   44631: out<=1;
   44632: out<=0;
   44633: out<=1;
   44634: out<=1;
   44635: out<=0;
   44636: out<=0;
   44637: out<=0;
   44638: out<=0;
   44639: out<=0;
   44640: out<=0;
   44641: out<=0;
   44642: out<=1;
   44643: out<=1;
   44644: out<=0;
   44645: out<=1;
   44646: out<=0;
   44647: out<=1;
   44648: out<=0;
   44649: out<=1;
   44650: out<=1;
   44651: out<=0;
   44652: out<=0;
   44653: out<=0;
   44654: out<=0;
   44655: out<=0;
   44656: out<=1;
   44657: out<=1;
   44658: out<=0;
   44659: out<=0;
   44660: out<=1;
   44661: out<=0;
   44662: out<=1;
   44663: out<=0;
   44664: out<=1;
   44665: out<=0;
   44666: out<=0;
   44667: out<=1;
   44668: out<=1;
   44669: out<=1;
   44670: out<=1;
   44671: out<=1;
   44672: out<=1;
   44673: out<=1;
   44674: out<=0;
   44675: out<=0;
   44676: out<=1;
   44677: out<=0;
   44678: out<=1;
   44679: out<=0;
   44680: out<=1;
   44681: out<=0;
   44682: out<=0;
   44683: out<=1;
   44684: out<=1;
   44685: out<=1;
   44686: out<=1;
   44687: out<=1;
   44688: out<=0;
   44689: out<=0;
   44690: out<=1;
   44691: out<=1;
   44692: out<=0;
   44693: out<=1;
   44694: out<=0;
   44695: out<=1;
   44696: out<=0;
   44697: out<=1;
   44698: out<=1;
   44699: out<=0;
   44700: out<=0;
   44701: out<=0;
   44702: out<=0;
   44703: out<=0;
   44704: out<=1;
   44705: out<=1;
   44706: out<=0;
   44707: out<=0;
   44708: out<=1;
   44709: out<=0;
   44710: out<=1;
   44711: out<=0;
   44712: out<=1;
   44713: out<=0;
   44714: out<=0;
   44715: out<=1;
   44716: out<=1;
   44717: out<=1;
   44718: out<=1;
   44719: out<=1;
   44720: out<=0;
   44721: out<=0;
   44722: out<=1;
   44723: out<=1;
   44724: out<=0;
   44725: out<=1;
   44726: out<=0;
   44727: out<=1;
   44728: out<=0;
   44729: out<=1;
   44730: out<=1;
   44731: out<=0;
   44732: out<=0;
   44733: out<=0;
   44734: out<=0;
   44735: out<=0;
   44736: out<=1;
   44737: out<=1;
   44738: out<=0;
   44739: out<=0;
   44740: out<=1;
   44741: out<=0;
   44742: out<=1;
   44743: out<=0;
   44744: out<=1;
   44745: out<=0;
   44746: out<=0;
   44747: out<=1;
   44748: out<=1;
   44749: out<=1;
   44750: out<=1;
   44751: out<=1;
   44752: out<=1;
   44753: out<=1;
   44754: out<=0;
   44755: out<=0;
   44756: out<=1;
   44757: out<=0;
   44758: out<=1;
   44759: out<=0;
   44760: out<=1;
   44761: out<=0;
   44762: out<=0;
   44763: out<=1;
   44764: out<=1;
   44765: out<=1;
   44766: out<=1;
   44767: out<=1;
   44768: out<=0;
   44769: out<=0;
   44770: out<=1;
   44771: out<=1;
   44772: out<=0;
   44773: out<=1;
   44774: out<=0;
   44775: out<=1;
   44776: out<=0;
   44777: out<=1;
   44778: out<=1;
   44779: out<=0;
   44780: out<=0;
   44781: out<=0;
   44782: out<=0;
   44783: out<=0;
   44784: out<=0;
   44785: out<=0;
   44786: out<=1;
   44787: out<=1;
   44788: out<=0;
   44789: out<=1;
   44790: out<=0;
   44791: out<=1;
   44792: out<=0;
   44793: out<=1;
   44794: out<=1;
   44795: out<=0;
   44796: out<=0;
   44797: out<=0;
   44798: out<=0;
   44799: out<=0;
   44800: out<=1;
   44801: out<=0;
   44802: out<=1;
   44803: out<=0;
   44804: out<=0;
   44805: out<=0;
   44806: out<=1;
   44807: out<=1;
   44808: out<=0;
   44809: out<=0;
   44810: out<=0;
   44811: out<=0;
   44812: out<=1;
   44813: out<=0;
   44814: out<=0;
   44815: out<=1;
   44816: out<=0;
   44817: out<=1;
   44818: out<=0;
   44819: out<=1;
   44820: out<=1;
   44821: out<=1;
   44822: out<=0;
   44823: out<=0;
   44824: out<=1;
   44825: out<=1;
   44826: out<=1;
   44827: out<=1;
   44828: out<=0;
   44829: out<=1;
   44830: out<=1;
   44831: out<=0;
   44832: out<=0;
   44833: out<=1;
   44834: out<=0;
   44835: out<=1;
   44836: out<=1;
   44837: out<=1;
   44838: out<=0;
   44839: out<=0;
   44840: out<=1;
   44841: out<=1;
   44842: out<=1;
   44843: out<=1;
   44844: out<=0;
   44845: out<=1;
   44846: out<=1;
   44847: out<=0;
   44848: out<=1;
   44849: out<=0;
   44850: out<=1;
   44851: out<=0;
   44852: out<=0;
   44853: out<=0;
   44854: out<=1;
   44855: out<=1;
   44856: out<=0;
   44857: out<=0;
   44858: out<=0;
   44859: out<=0;
   44860: out<=1;
   44861: out<=0;
   44862: out<=0;
   44863: out<=1;
   44864: out<=1;
   44865: out<=0;
   44866: out<=1;
   44867: out<=0;
   44868: out<=0;
   44869: out<=0;
   44870: out<=1;
   44871: out<=1;
   44872: out<=0;
   44873: out<=0;
   44874: out<=0;
   44875: out<=0;
   44876: out<=1;
   44877: out<=0;
   44878: out<=0;
   44879: out<=1;
   44880: out<=1;
   44881: out<=0;
   44882: out<=1;
   44883: out<=0;
   44884: out<=0;
   44885: out<=0;
   44886: out<=1;
   44887: out<=1;
   44888: out<=0;
   44889: out<=0;
   44890: out<=0;
   44891: out<=0;
   44892: out<=1;
   44893: out<=0;
   44894: out<=0;
   44895: out<=1;
   44896: out<=1;
   44897: out<=0;
   44898: out<=1;
   44899: out<=0;
   44900: out<=0;
   44901: out<=0;
   44902: out<=1;
   44903: out<=1;
   44904: out<=0;
   44905: out<=0;
   44906: out<=0;
   44907: out<=0;
   44908: out<=1;
   44909: out<=0;
   44910: out<=0;
   44911: out<=1;
   44912: out<=1;
   44913: out<=0;
   44914: out<=1;
   44915: out<=0;
   44916: out<=0;
   44917: out<=0;
   44918: out<=1;
   44919: out<=1;
   44920: out<=0;
   44921: out<=0;
   44922: out<=0;
   44923: out<=0;
   44924: out<=1;
   44925: out<=0;
   44926: out<=0;
   44927: out<=1;
   44928: out<=1;
   44929: out<=0;
   44930: out<=1;
   44931: out<=0;
   44932: out<=0;
   44933: out<=0;
   44934: out<=1;
   44935: out<=1;
   44936: out<=0;
   44937: out<=0;
   44938: out<=0;
   44939: out<=0;
   44940: out<=1;
   44941: out<=0;
   44942: out<=0;
   44943: out<=1;
   44944: out<=1;
   44945: out<=0;
   44946: out<=1;
   44947: out<=0;
   44948: out<=0;
   44949: out<=0;
   44950: out<=1;
   44951: out<=1;
   44952: out<=0;
   44953: out<=0;
   44954: out<=0;
   44955: out<=0;
   44956: out<=1;
   44957: out<=0;
   44958: out<=0;
   44959: out<=1;
   44960: out<=0;
   44961: out<=1;
   44962: out<=0;
   44963: out<=1;
   44964: out<=1;
   44965: out<=1;
   44966: out<=0;
   44967: out<=0;
   44968: out<=1;
   44969: out<=1;
   44970: out<=1;
   44971: out<=1;
   44972: out<=0;
   44973: out<=1;
   44974: out<=1;
   44975: out<=0;
   44976: out<=0;
   44977: out<=1;
   44978: out<=0;
   44979: out<=1;
   44980: out<=1;
   44981: out<=1;
   44982: out<=0;
   44983: out<=0;
   44984: out<=1;
   44985: out<=1;
   44986: out<=1;
   44987: out<=1;
   44988: out<=0;
   44989: out<=1;
   44990: out<=1;
   44991: out<=0;
   44992: out<=1;
   44993: out<=0;
   44994: out<=1;
   44995: out<=0;
   44996: out<=0;
   44997: out<=0;
   44998: out<=1;
   44999: out<=1;
   45000: out<=0;
   45001: out<=0;
   45002: out<=0;
   45003: out<=0;
   45004: out<=1;
   45005: out<=0;
   45006: out<=0;
   45007: out<=1;
   45008: out<=0;
   45009: out<=1;
   45010: out<=0;
   45011: out<=1;
   45012: out<=1;
   45013: out<=1;
   45014: out<=0;
   45015: out<=0;
   45016: out<=1;
   45017: out<=1;
   45018: out<=1;
   45019: out<=1;
   45020: out<=0;
   45021: out<=1;
   45022: out<=1;
   45023: out<=0;
   45024: out<=1;
   45025: out<=0;
   45026: out<=1;
   45027: out<=0;
   45028: out<=0;
   45029: out<=0;
   45030: out<=1;
   45031: out<=1;
   45032: out<=0;
   45033: out<=0;
   45034: out<=0;
   45035: out<=0;
   45036: out<=1;
   45037: out<=0;
   45038: out<=0;
   45039: out<=1;
   45040: out<=0;
   45041: out<=1;
   45042: out<=0;
   45043: out<=1;
   45044: out<=1;
   45045: out<=1;
   45046: out<=0;
   45047: out<=0;
   45048: out<=1;
   45049: out<=1;
   45050: out<=1;
   45051: out<=1;
   45052: out<=0;
   45053: out<=1;
   45054: out<=1;
   45055: out<=0;
   45056: out<=1;
   45057: out<=1;
   45058: out<=0;
   45059: out<=0;
   45060: out<=0;
   45061: out<=1;
   45062: out<=0;
   45063: out<=1;
   45064: out<=1;
   45065: out<=0;
   45066: out<=0;
   45067: out<=1;
   45068: out<=0;
   45069: out<=0;
   45070: out<=0;
   45071: out<=0;
   45072: out<=1;
   45073: out<=1;
   45074: out<=0;
   45075: out<=0;
   45076: out<=0;
   45077: out<=1;
   45078: out<=0;
   45079: out<=1;
   45080: out<=1;
   45081: out<=0;
   45082: out<=0;
   45083: out<=1;
   45084: out<=0;
   45085: out<=0;
   45086: out<=0;
   45087: out<=0;
   45088: out<=0;
   45089: out<=0;
   45090: out<=1;
   45091: out<=1;
   45092: out<=1;
   45093: out<=0;
   45094: out<=1;
   45095: out<=0;
   45096: out<=0;
   45097: out<=1;
   45098: out<=1;
   45099: out<=0;
   45100: out<=1;
   45101: out<=1;
   45102: out<=1;
   45103: out<=1;
   45104: out<=0;
   45105: out<=0;
   45106: out<=1;
   45107: out<=1;
   45108: out<=1;
   45109: out<=0;
   45110: out<=1;
   45111: out<=0;
   45112: out<=0;
   45113: out<=1;
   45114: out<=1;
   45115: out<=0;
   45116: out<=1;
   45117: out<=1;
   45118: out<=1;
   45119: out<=1;
   45120: out<=0;
   45121: out<=0;
   45122: out<=1;
   45123: out<=1;
   45124: out<=1;
   45125: out<=0;
   45126: out<=1;
   45127: out<=0;
   45128: out<=0;
   45129: out<=1;
   45130: out<=1;
   45131: out<=0;
   45132: out<=1;
   45133: out<=1;
   45134: out<=1;
   45135: out<=1;
   45136: out<=1;
   45137: out<=1;
   45138: out<=0;
   45139: out<=0;
   45140: out<=0;
   45141: out<=1;
   45142: out<=0;
   45143: out<=1;
   45144: out<=1;
   45145: out<=0;
   45146: out<=0;
   45147: out<=1;
   45148: out<=0;
   45149: out<=0;
   45150: out<=0;
   45151: out<=0;
   45152: out<=0;
   45153: out<=0;
   45154: out<=1;
   45155: out<=1;
   45156: out<=1;
   45157: out<=0;
   45158: out<=1;
   45159: out<=0;
   45160: out<=0;
   45161: out<=1;
   45162: out<=1;
   45163: out<=0;
   45164: out<=1;
   45165: out<=1;
   45166: out<=1;
   45167: out<=1;
   45168: out<=1;
   45169: out<=1;
   45170: out<=0;
   45171: out<=0;
   45172: out<=0;
   45173: out<=1;
   45174: out<=0;
   45175: out<=1;
   45176: out<=1;
   45177: out<=0;
   45178: out<=0;
   45179: out<=1;
   45180: out<=0;
   45181: out<=0;
   45182: out<=0;
   45183: out<=0;
   45184: out<=0;
   45185: out<=0;
   45186: out<=1;
   45187: out<=1;
   45188: out<=1;
   45189: out<=0;
   45190: out<=1;
   45191: out<=0;
   45192: out<=0;
   45193: out<=1;
   45194: out<=1;
   45195: out<=0;
   45196: out<=1;
   45197: out<=1;
   45198: out<=1;
   45199: out<=1;
   45200: out<=1;
   45201: out<=1;
   45202: out<=0;
   45203: out<=0;
   45204: out<=0;
   45205: out<=1;
   45206: out<=0;
   45207: out<=1;
   45208: out<=1;
   45209: out<=0;
   45210: out<=0;
   45211: out<=1;
   45212: out<=0;
   45213: out<=0;
   45214: out<=0;
   45215: out<=0;
   45216: out<=1;
   45217: out<=1;
   45218: out<=0;
   45219: out<=0;
   45220: out<=0;
   45221: out<=1;
   45222: out<=0;
   45223: out<=1;
   45224: out<=1;
   45225: out<=0;
   45226: out<=0;
   45227: out<=1;
   45228: out<=0;
   45229: out<=0;
   45230: out<=0;
   45231: out<=0;
   45232: out<=0;
   45233: out<=0;
   45234: out<=1;
   45235: out<=1;
   45236: out<=1;
   45237: out<=0;
   45238: out<=1;
   45239: out<=0;
   45240: out<=0;
   45241: out<=1;
   45242: out<=1;
   45243: out<=0;
   45244: out<=1;
   45245: out<=1;
   45246: out<=1;
   45247: out<=1;
   45248: out<=1;
   45249: out<=1;
   45250: out<=0;
   45251: out<=0;
   45252: out<=0;
   45253: out<=1;
   45254: out<=0;
   45255: out<=1;
   45256: out<=1;
   45257: out<=0;
   45258: out<=0;
   45259: out<=1;
   45260: out<=0;
   45261: out<=0;
   45262: out<=0;
   45263: out<=0;
   45264: out<=1;
   45265: out<=1;
   45266: out<=0;
   45267: out<=0;
   45268: out<=0;
   45269: out<=1;
   45270: out<=0;
   45271: out<=1;
   45272: out<=1;
   45273: out<=0;
   45274: out<=0;
   45275: out<=1;
   45276: out<=0;
   45277: out<=0;
   45278: out<=0;
   45279: out<=0;
   45280: out<=1;
   45281: out<=1;
   45282: out<=0;
   45283: out<=0;
   45284: out<=0;
   45285: out<=1;
   45286: out<=0;
   45287: out<=1;
   45288: out<=1;
   45289: out<=0;
   45290: out<=0;
   45291: out<=1;
   45292: out<=0;
   45293: out<=0;
   45294: out<=0;
   45295: out<=0;
   45296: out<=1;
   45297: out<=1;
   45298: out<=0;
   45299: out<=0;
   45300: out<=0;
   45301: out<=1;
   45302: out<=0;
   45303: out<=1;
   45304: out<=1;
   45305: out<=0;
   45306: out<=0;
   45307: out<=1;
   45308: out<=0;
   45309: out<=0;
   45310: out<=0;
   45311: out<=0;
   45312: out<=1;
   45313: out<=0;
   45314: out<=1;
   45315: out<=0;
   45316: out<=1;
   45317: out<=1;
   45318: out<=0;
   45319: out<=0;
   45320: out<=0;
   45321: out<=0;
   45322: out<=0;
   45323: out<=0;
   45324: out<=0;
   45325: out<=1;
   45326: out<=1;
   45327: out<=0;
   45328: out<=0;
   45329: out<=1;
   45330: out<=0;
   45331: out<=1;
   45332: out<=0;
   45333: out<=0;
   45334: out<=1;
   45335: out<=1;
   45336: out<=1;
   45337: out<=1;
   45338: out<=1;
   45339: out<=1;
   45340: out<=1;
   45341: out<=0;
   45342: out<=0;
   45343: out<=1;
   45344: out<=1;
   45345: out<=0;
   45346: out<=1;
   45347: out<=0;
   45348: out<=1;
   45349: out<=1;
   45350: out<=0;
   45351: out<=0;
   45352: out<=0;
   45353: out<=0;
   45354: out<=0;
   45355: out<=0;
   45356: out<=0;
   45357: out<=1;
   45358: out<=1;
   45359: out<=0;
   45360: out<=0;
   45361: out<=1;
   45362: out<=0;
   45363: out<=1;
   45364: out<=0;
   45365: out<=0;
   45366: out<=1;
   45367: out<=1;
   45368: out<=1;
   45369: out<=1;
   45370: out<=1;
   45371: out<=1;
   45372: out<=1;
   45373: out<=0;
   45374: out<=0;
   45375: out<=1;
   45376: out<=0;
   45377: out<=1;
   45378: out<=0;
   45379: out<=1;
   45380: out<=0;
   45381: out<=0;
   45382: out<=1;
   45383: out<=1;
   45384: out<=1;
   45385: out<=1;
   45386: out<=1;
   45387: out<=1;
   45388: out<=1;
   45389: out<=0;
   45390: out<=0;
   45391: out<=1;
   45392: out<=0;
   45393: out<=1;
   45394: out<=0;
   45395: out<=1;
   45396: out<=0;
   45397: out<=0;
   45398: out<=1;
   45399: out<=1;
   45400: out<=1;
   45401: out<=1;
   45402: out<=1;
   45403: out<=1;
   45404: out<=1;
   45405: out<=0;
   45406: out<=0;
   45407: out<=1;
   45408: out<=1;
   45409: out<=0;
   45410: out<=1;
   45411: out<=0;
   45412: out<=1;
   45413: out<=1;
   45414: out<=0;
   45415: out<=0;
   45416: out<=0;
   45417: out<=0;
   45418: out<=0;
   45419: out<=0;
   45420: out<=0;
   45421: out<=1;
   45422: out<=1;
   45423: out<=0;
   45424: out<=1;
   45425: out<=0;
   45426: out<=1;
   45427: out<=0;
   45428: out<=1;
   45429: out<=1;
   45430: out<=0;
   45431: out<=0;
   45432: out<=0;
   45433: out<=0;
   45434: out<=0;
   45435: out<=0;
   45436: out<=0;
   45437: out<=1;
   45438: out<=1;
   45439: out<=0;
   45440: out<=0;
   45441: out<=1;
   45442: out<=0;
   45443: out<=1;
   45444: out<=0;
   45445: out<=0;
   45446: out<=1;
   45447: out<=1;
   45448: out<=1;
   45449: out<=1;
   45450: out<=1;
   45451: out<=1;
   45452: out<=1;
   45453: out<=0;
   45454: out<=0;
   45455: out<=1;
   45456: out<=0;
   45457: out<=1;
   45458: out<=0;
   45459: out<=1;
   45460: out<=0;
   45461: out<=0;
   45462: out<=1;
   45463: out<=1;
   45464: out<=1;
   45465: out<=1;
   45466: out<=1;
   45467: out<=1;
   45468: out<=1;
   45469: out<=0;
   45470: out<=0;
   45471: out<=1;
   45472: out<=0;
   45473: out<=1;
   45474: out<=0;
   45475: out<=1;
   45476: out<=0;
   45477: out<=0;
   45478: out<=1;
   45479: out<=1;
   45480: out<=1;
   45481: out<=1;
   45482: out<=1;
   45483: out<=1;
   45484: out<=1;
   45485: out<=0;
   45486: out<=0;
   45487: out<=1;
   45488: out<=0;
   45489: out<=1;
   45490: out<=0;
   45491: out<=1;
   45492: out<=0;
   45493: out<=0;
   45494: out<=1;
   45495: out<=1;
   45496: out<=1;
   45497: out<=1;
   45498: out<=1;
   45499: out<=1;
   45500: out<=1;
   45501: out<=0;
   45502: out<=0;
   45503: out<=1;
   45504: out<=1;
   45505: out<=0;
   45506: out<=1;
   45507: out<=0;
   45508: out<=1;
   45509: out<=1;
   45510: out<=0;
   45511: out<=0;
   45512: out<=0;
   45513: out<=0;
   45514: out<=0;
   45515: out<=0;
   45516: out<=0;
   45517: out<=1;
   45518: out<=1;
   45519: out<=0;
   45520: out<=0;
   45521: out<=1;
   45522: out<=0;
   45523: out<=1;
   45524: out<=0;
   45525: out<=0;
   45526: out<=1;
   45527: out<=1;
   45528: out<=1;
   45529: out<=1;
   45530: out<=1;
   45531: out<=1;
   45532: out<=1;
   45533: out<=0;
   45534: out<=0;
   45535: out<=1;
   45536: out<=0;
   45537: out<=1;
   45538: out<=0;
   45539: out<=1;
   45540: out<=0;
   45541: out<=0;
   45542: out<=1;
   45543: out<=1;
   45544: out<=1;
   45545: out<=1;
   45546: out<=1;
   45547: out<=1;
   45548: out<=1;
   45549: out<=0;
   45550: out<=0;
   45551: out<=1;
   45552: out<=1;
   45553: out<=0;
   45554: out<=1;
   45555: out<=0;
   45556: out<=1;
   45557: out<=1;
   45558: out<=0;
   45559: out<=0;
   45560: out<=0;
   45561: out<=0;
   45562: out<=0;
   45563: out<=0;
   45564: out<=0;
   45565: out<=1;
   45566: out<=1;
   45567: out<=0;
   45568: out<=1;
   45569: out<=0;
   45570: out<=0;
   45571: out<=1;
   45572: out<=1;
   45573: out<=1;
   45574: out<=1;
   45575: out<=1;
   45576: out<=1;
   45577: out<=1;
   45578: out<=0;
   45579: out<=0;
   45580: out<=1;
   45581: out<=0;
   45582: out<=1;
   45583: out<=0;
   45584: out<=0;
   45585: out<=1;
   45586: out<=1;
   45587: out<=0;
   45588: out<=0;
   45589: out<=0;
   45590: out<=0;
   45591: out<=0;
   45592: out<=0;
   45593: out<=0;
   45594: out<=1;
   45595: out<=1;
   45596: out<=0;
   45597: out<=1;
   45598: out<=0;
   45599: out<=1;
   45600: out<=0;
   45601: out<=1;
   45602: out<=1;
   45603: out<=0;
   45604: out<=0;
   45605: out<=0;
   45606: out<=0;
   45607: out<=0;
   45608: out<=0;
   45609: out<=0;
   45610: out<=1;
   45611: out<=1;
   45612: out<=0;
   45613: out<=1;
   45614: out<=0;
   45615: out<=1;
   45616: out<=1;
   45617: out<=0;
   45618: out<=0;
   45619: out<=1;
   45620: out<=1;
   45621: out<=1;
   45622: out<=1;
   45623: out<=1;
   45624: out<=1;
   45625: out<=1;
   45626: out<=0;
   45627: out<=0;
   45628: out<=1;
   45629: out<=0;
   45630: out<=1;
   45631: out<=0;
   45632: out<=0;
   45633: out<=1;
   45634: out<=1;
   45635: out<=0;
   45636: out<=0;
   45637: out<=0;
   45638: out<=0;
   45639: out<=0;
   45640: out<=0;
   45641: out<=0;
   45642: out<=1;
   45643: out<=1;
   45644: out<=0;
   45645: out<=1;
   45646: out<=0;
   45647: out<=1;
   45648: out<=0;
   45649: out<=1;
   45650: out<=1;
   45651: out<=0;
   45652: out<=0;
   45653: out<=0;
   45654: out<=0;
   45655: out<=0;
   45656: out<=0;
   45657: out<=0;
   45658: out<=1;
   45659: out<=1;
   45660: out<=0;
   45661: out<=1;
   45662: out<=0;
   45663: out<=1;
   45664: out<=0;
   45665: out<=1;
   45666: out<=1;
   45667: out<=0;
   45668: out<=0;
   45669: out<=0;
   45670: out<=0;
   45671: out<=0;
   45672: out<=0;
   45673: out<=0;
   45674: out<=1;
   45675: out<=1;
   45676: out<=0;
   45677: out<=1;
   45678: out<=0;
   45679: out<=1;
   45680: out<=0;
   45681: out<=1;
   45682: out<=1;
   45683: out<=0;
   45684: out<=0;
   45685: out<=0;
   45686: out<=0;
   45687: out<=0;
   45688: out<=0;
   45689: out<=0;
   45690: out<=1;
   45691: out<=1;
   45692: out<=0;
   45693: out<=1;
   45694: out<=0;
   45695: out<=1;
   45696: out<=0;
   45697: out<=1;
   45698: out<=1;
   45699: out<=0;
   45700: out<=0;
   45701: out<=0;
   45702: out<=0;
   45703: out<=0;
   45704: out<=0;
   45705: out<=0;
   45706: out<=1;
   45707: out<=1;
   45708: out<=0;
   45709: out<=1;
   45710: out<=0;
   45711: out<=1;
   45712: out<=0;
   45713: out<=1;
   45714: out<=1;
   45715: out<=0;
   45716: out<=0;
   45717: out<=0;
   45718: out<=0;
   45719: out<=0;
   45720: out<=0;
   45721: out<=0;
   45722: out<=1;
   45723: out<=1;
   45724: out<=0;
   45725: out<=1;
   45726: out<=0;
   45727: out<=1;
   45728: out<=1;
   45729: out<=0;
   45730: out<=0;
   45731: out<=1;
   45732: out<=1;
   45733: out<=1;
   45734: out<=1;
   45735: out<=1;
   45736: out<=1;
   45737: out<=1;
   45738: out<=0;
   45739: out<=0;
   45740: out<=1;
   45741: out<=0;
   45742: out<=1;
   45743: out<=0;
   45744: out<=1;
   45745: out<=0;
   45746: out<=0;
   45747: out<=1;
   45748: out<=1;
   45749: out<=1;
   45750: out<=1;
   45751: out<=1;
   45752: out<=1;
   45753: out<=1;
   45754: out<=0;
   45755: out<=0;
   45756: out<=1;
   45757: out<=0;
   45758: out<=1;
   45759: out<=0;
   45760: out<=1;
   45761: out<=0;
   45762: out<=0;
   45763: out<=1;
   45764: out<=1;
   45765: out<=1;
   45766: out<=1;
   45767: out<=1;
   45768: out<=1;
   45769: out<=1;
   45770: out<=0;
   45771: out<=0;
   45772: out<=1;
   45773: out<=0;
   45774: out<=1;
   45775: out<=0;
   45776: out<=0;
   45777: out<=1;
   45778: out<=1;
   45779: out<=0;
   45780: out<=0;
   45781: out<=0;
   45782: out<=0;
   45783: out<=0;
   45784: out<=0;
   45785: out<=0;
   45786: out<=1;
   45787: out<=1;
   45788: out<=0;
   45789: out<=1;
   45790: out<=0;
   45791: out<=1;
   45792: out<=1;
   45793: out<=0;
   45794: out<=0;
   45795: out<=1;
   45796: out<=1;
   45797: out<=1;
   45798: out<=1;
   45799: out<=1;
   45800: out<=1;
   45801: out<=1;
   45802: out<=0;
   45803: out<=0;
   45804: out<=1;
   45805: out<=0;
   45806: out<=1;
   45807: out<=0;
   45808: out<=0;
   45809: out<=1;
   45810: out<=1;
   45811: out<=0;
   45812: out<=0;
   45813: out<=0;
   45814: out<=0;
   45815: out<=0;
   45816: out<=0;
   45817: out<=0;
   45818: out<=1;
   45819: out<=1;
   45820: out<=0;
   45821: out<=1;
   45822: out<=0;
   45823: out<=1;
   45824: out<=1;
   45825: out<=1;
   45826: out<=1;
   45827: out<=1;
   45828: out<=0;
   45829: out<=1;
   45830: out<=1;
   45831: out<=0;
   45832: out<=0;
   45833: out<=1;
   45834: out<=0;
   45835: out<=1;
   45836: out<=1;
   45837: out<=1;
   45838: out<=0;
   45839: out<=0;
   45840: out<=1;
   45841: out<=1;
   45842: out<=1;
   45843: out<=1;
   45844: out<=0;
   45845: out<=1;
   45846: out<=1;
   45847: out<=0;
   45848: out<=0;
   45849: out<=1;
   45850: out<=0;
   45851: out<=1;
   45852: out<=1;
   45853: out<=1;
   45854: out<=0;
   45855: out<=0;
   45856: out<=1;
   45857: out<=1;
   45858: out<=1;
   45859: out<=1;
   45860: out<=0;
   45861: out<=1;
   45862: out<=1;
   45863: out<=0;
   45864: out<=0;
   45865: out<=1;
   45866: out<=0;
   45867: out<=1;
   45868: out<=1;
   45869: out<=1;
   45870: out<=0;
   45871: out<=0;
   45872: out<=1;
   45873: out<=1;
   45874: out<=1;
   45875: out<=1;
   45876: out<=0;
   45877: out<=1;
   45878: out<=1;
   45879: out<=0;
   45880: out<=0;
   45881: out<=1;
   45882: out<=0;
   45883: out<=1;
   45884: out<=1;
   45885: out<=1;
   45886: out<=0;
   45887: out<=0;
   45888: out<=0;
   45889: out<=0;
   45890: out<=0;
   45891: out<=0;
   45892: out<=1;
   45893: out<=0;
   45894: out<=0;
   45895: out<=1;
   45896: out<=1;
   45897: out<=0;
   45898: out<=1;
   45899: out<=0;
   45900: out<=0;
   45901: out<=0;
   45902: out<=1;
   45903: out<=1;
   45904: out<=1;
   45905: out<=1;
   45906: out<=1;
   45907: out<=1;
   45908: out<=0;
   45909: out<=1;
   45910: out<=1;
   45911: out<=0;
   45912: out<=0;
   45913: out<=1;
   45914: out<=0;
   45915: out<=1;
   45916: out<=1;
   45917: out<=1;
   45918: out<=0;
   45919: out<=0;
   45920: out<=1;
   45921: out<=1;
   45922: out<=1;
   45923: out<=1;
   45924: out<=0;
   45925: out<=1;
   45926: out<=1;
   45927: out<=0;
   45928: out<=0;
   45929: out<=1;
   45930: out<=0;
   45931: out<=1;
   45932: out<=1;
   45933: out<=1;
   45934: out<=0;
   45935: out<=0;
   45936: out<=0;
   45937: out<=0;
   45938: out<=0;
   45939: out<=0;
   45940: out<=1;
   45941: out<=0;
   45942: out<=0;
   45943: out<=1;
   45944: out<=1;
   45945: out<=0;
   45946: out<=1;
   45947: out<=0;
   45948: out<=0;
   45949: out<=0;
   45950: out<=1;
   45951: out<=1;
   45952: out<=0;
   45953: out<=0;
   45954: out<=0;
   45955: out<=0;
   45956: out<=1;
   45957: out<=0;
   45958: out<=0;
   45959: out<=1;
   45960: out<=1;
   45961: out<=0;
   45962: out<=1;
   45963: out<=0;
   45964: out<=0;
   45965: out<=0;
   45966: out<=1;
   45967: out<=1;
   45968: out<=1;
   45969: out<=1;
   45970: out<=1;
   45971: out<=1;
   45972: out<=0;
   45973: out<=1;
   45974: out<=1;
   45975: out<=0;
   45976: out<=0;
   45977: out<=1;
   45978: out<=0;
   45979: out<=1;
   45980: out<=1;
   45981: out<=1;
   45982: out<=0;
   45983: out<=0;
   45984: out<=0;
   45985: out<=0;
   45986: out<=0;
   45987: out<=0;
   45988: out<=1;
   45989: out<=0;
   45990: out<=0;
   45991: out<=1;
   45992: out<=1;
   45993: out<=0;
   45994: out<=1;
   45995: out<=0;
   45996: out<=0;
   45997: out<=0;
   45998: out<=1;
   45999: out<=1;
   46000: out<=1;
   46001: out<=1;
   46002: out<=1;
   46003: out<=1;
   46004: out<=0;
   46005: out<=1;
   46006: out<=1;
   46007: out<=0;
   46008: out<=0;
   46009: out<=1;
   46010: out<=0;
   46011: out<=1;
   46012: out<=1;
   46013: out<=1;
   46014: out<=0;
   46015: out<=0;
   46016: out<=1;
   46017: out<=1;
   46018: out<=1;
   46019: out<=1;
   46020: out<=0;
   46021: out<=1;
   46022: out<=1;
   46023: out<=0;
   46024: out<=0;
   46025: out<=1;
   46026: out<=0;
   46027: out<=1;
   46028: out<=1;
   46029: out<=1;
   46030: out<=0;
   46031: out<=0;
   46032: out<=1;
   46033: out<=1;
   46034: out<=1;
   46035: out<=1;
   46036: out<=0;
   46037: out<=1;
   46038: out<=1;
   46039: out<=0;
   46040: out<=0;
   46041: out<=1;
   46042: out<=0;
   46043: out<=1;
   46044: out<=1;
   46045: out<=1;
   46046: out<=0;
   46047: out<=0;
   46048: out<=0;
   46049: out<=0;
   46050: out<=0;
   46051: out<=0;
   46052: out<=1;
   46053: out<=0;
   46054: out<=0;
   46055: out<=1;
   46056: out<=1;
   46057: out<=0;
   46058: out<=1;
   46059: out<=0;
   46060: out<=0;
   46061: out<=0;
   46062: out<=1;
   46063: out<=1;
   46064: out<=0;
   46065: out<=0;
   46066: out<=0;
   46067: out<=0;
   46068: out<=1;
   46069: out<=0;
   46070: out<=0;
   46071: out<=1;
   46072: out<=1;
   46073: out<=0;
   46074: out<=1;
   46075: out<=0;
   46076: out<=0;
   46077: out<=0;
   46078: out<=1;
   46079: out<=1;
   46080: out<=1;
   46081: out<=0;
   46082: out<=1;
   46083: out<=0;
   46084: out<=0;
   46085: out<=0;
   46086: out<=1;
   46087: out<=1;
   46088: out<=1;
   46089: out<=1;
   46090: out<=1;
   46091: out<=1;
   46092: out<=0;
   46093: out<=1;
   46094: out<=1;
   46095: out<=0;
   46096: out<=1;
   46097: out<=0;
   46098: out<=1;
   46099: out<=0;
   46100: out<=0;
   46101: out<=0;
   46102: out<=1;
   46103: out<=1;
   46104: out<=1;
   46105: out<=1;
   46106: out<=1;
   46107: out<=1;
   46108: out<=0;
   46109: out<=1;
   46110: out<=1;
   46111: out<=0;
   46112: out<=0;
   46113: out<=1;
   46114: out<=0;
   46115: out<=1;
   46116: out<=1;
   46117: out<=1;
   46118: out<=0;
   46119: out<=0;
   46120: out<=0;
   46121: out<=0;
   46122: out<=0;
   46123: out<=0;
   46124: out<=1;
   46125: out<=0;
   46126: out<=0;
   46127: out<=1;
   46128: out<=0;
   46129: out<=1;
   46130: out<=0;
   46131: out<=1;
   46132: out<=1;
   46133: out<=1;
   46134: out<=0;
   46135: out<=0;
   46136: out<=0;
   46137: out<=0;
   46138: out<=0;
   46139: out<=0;
   46140: out<=1;
   46141: out<=0;
   46142: out<=0;
   46143: out<=1;
   46144: out<=0;
   46145: out<=1;
   46146: out<=0;
   46147: out<=1;
   46148: out<=1;
   46149: out<=1;
   46150: out<=0;
   46151: out<=0;
   46152: out<=0;
   46153: out<=0;
   46154: out<=0;
   46155: out<=0;
   46156: out<=1;
   46157: out<=0;
   46158: out<=0;
   46159: out<=1;
   46160: out<=1;
   46161: out<=0;
   46162: out<=1;
   46163: out<=0;
   46164: out<=0;
   46165: out<=0;
   46166: out<=1;
   46167: out<=1;
   46168: out<=1;
   46169: out<=1;
   46170: out<=1;
   46171: out<=1;
   46172: out<=0;
   46173: out<=1;
   46174: out<=1;
   46175: out<=0;
   46176: out<=0;
   46177: out<=1;
   46178: out<=0;
   46179: out<=1;
   46180: out<=1;
   46181: out<=1;
   46182: out<=0;
   46183: out<=0;
   46184: out<=0;
   46185: out<=0;
   46186: out<=0;
   46187: out<=0;
   46188: out<=1;
   46189: out<=0;
   46190: out<=0;
   46191: out<=1;
   46192: out<=1;
   46193: out<=0;
   46194: out<=1;
   46195: out<=0;
   46196: out<=0;
   46197: out<=0;
   46198: out<=1;
   46199: out<=1;
   46200: out<=1;
   46201: out<=1;
   46202: out<=1;
   46203: out<=1;
   46204: out<=0;
   46205: out<=1;
   46206: out<=1;
   46207: out<=0;
   46208: out<=0;
   46209: out<=1;
   46210: out<=0;
   46211: out<=1;
   46212: out<=1;
   46213: out<=1;
   46214: out<=0;
   46215: out<=0;
   46216: out<=0;
   46217: out<=0;
   46218: out<=0;
   46219: out<=0;
   46220: out<=1;
   46221: out<=0;
   46222: out<=0;
   46223: out<=1;
   46224: out<=1;
   46225: out<=0;
   46226: out<=1;
   46227: out<=0;
   46228: out<=0;
   46229: out<=0;
   46230: out<=1;
   46231: out<=1;
   46232: out<=1;
   46233: out<=1;
   46234: out<=1;
   46235: out<=1;
   46236: out<=0;
   46237: out<=1;
   46238: out<=1;
   46239: out<=0;
   46240: out<=1;
   46241: out<=0;
   46242: out<=1;
   46243: out<=0;
   46244: out<=0;
   46245: out<=0;
   46246: out<=1;
   46247: out<=1;
   46248: out<=1;
   46249: out<=1;
   46250: out<=1;
   46251: out<=1;
   46252: out<=0;
   46253: out<=1;
   46254: out<=1;
   46255: out<=0;
   46256: out<=0;
   46257: out<=1;
   46258: out<=0;
   46259: out<=1;
   46260: out<=1;
   46261: out<=1;
   46262: out<=0;
   46263: out<=0;
   46264: out<=0;
   46265: out<=0;
   46266: out<=0;
   46267: out<=0;
   46268: out<=1;
   46269: out<=0;
   46270: out<=0;
   46271: out<=1;
   46272: out<=1;
   46273: out<=0;
   46274: out<=1;
   46275: out<=0;
   46276: out<=0;
   46277: out<=0;
   46278: out<=1;
   46279: out<=1;
   46280: out<=1;
   46281: out<=1;
   46282: out<=1;
   46283: out<=1;
   46284: out<=0;
   46285: out<=1;
   46286: out<=1;
   46287: out<=0;
   46288: out<=1;
   46289: out<=0;
   46290: out<=1;
   46291: out<=0;
   46292: out<=0;
   46293: out<=0;
   46294: out<=1;
   46295: out<=1;
   46296: out<=1;
   46297: out<=1;
   46298: out<=1;
   46299: out<=1;
   46300: out<=0;
   46301: out<=1;
   46302: out<=1;
   46303: out<=0;
   46304: out<=1;
   46305: out<=0;
   46306: out<=1;
   46307: out<=0;
   46308: out<=0;
   46309: out<=0;
   46310: out<=1;
   46311: out<=1;
   46312: out<=1;
   46313: out<=1;
   46314: out<=1;
   46315: out<=1;
   46316: out<=0;
   46317: out<=1;
   46318: out<=1;
   46319: out<=0;
   46320: out<=1;
   46321: out<=0;
   46322: out<=1;
   46323: out<=0;
   46324: out<=0;
   46325: out<=0;
   46326: out<=1;
   46327: out<=1;
   46328: out<=1;
   46329: out<=1;
   46330: out<=1;
   46331: out<=1;
   46332: out<=0;
   46333: out<=1;
   46334: out<=1;
   46335: out<=0;
   46336: out<=0;
   46337: out<=0;
   46338: out<=1;
   46339: out<=1;
   46340: out<=0;
   46341: out<=1;
   46342: out<=0;
   46343: out<=1;
   46344: out<=1;
   46345: out<=0;
   46346: out<=0;
   46347: out<=1;
   46348: out<=1;
   46349: out<=1;
   46350: out<=1;
   46351: out<=1;
   46352: out<=1;
   46353: out<=1;
   46354: out<=0;
   46355: out<=0;
   46356: out<=1;
   46357: out<=0;
   46358: out<=1;
   46359: out<=0;
   46360: out<=0;
   46361: out<=1;
   46362: out<=1;
   46363: out<=0;
   46364: out<=0;
   46365: out<=0;
   46366: out<=0;
   46367: out<=0;
   46368: out<=0;
   46369: out<=0;
   46370: out<=1;
   46371: out<=1;
   46372: out<=0;
   46373: out<=1;
   46374: out<=0;
   46375: out<=1;
   46376: out<=1;
   46377: out<=0;
   46378: out<=0;
   46379: out<=1;
   46380: out<=1;
   46381: out<=1;
   46382: out<=1;
   46383: out<=1;
   46384: out<=1;
   46385: out<=1;
   46386: out<=0;
   46387: out<=0;
   46388: out<=1;
   46389: out<=0;
   46390: out<=1;
   46391: out<=0;
   46392: out<=0;
   46393: out<=1;
   46394: out<=1;
   46395: out<=0;
   46396: out<=0;
   46397: out<=0;
   46398: out<=0;
   46399: out<=0;
   46400: out<=1;
   46401: out<=1;
   46402: out<=0;
   46403: out<=0;
   46404: out<=1;
   46405: out<=0;
   46406: out<=1;
   46407: out<=0;
   46408: out<=0;
   46409: out<=1;
   46410: out<=1;
   46411: out<=0;
   46412: out<=0;
   46413: out<=0;
   46414: out<=0;
   46415: out<=0;
   46416: out<=1;
   46417: out<=1;
   46418: out<=0;
   46419: out<=0;
   46420: out<=1;
   46421: out<=0;
   46422: out<=1;
   46423: out<=0;
   46424: out<=0;
   46425: out<=1;
   46426: out<=1;
   46427: out<=0;
   46428: out<=0;
   46429: out<=0;
   46430: out<=0;
   46431: out<=0;
   46432: out<=0;
   46433: out<=0;
   46434: out<=1;
   46435: out<=1;
   46436: out<=0;
   46437: out<=1;
   46438: out<=0;
   46439: out<=1;
   46440: out<=1;
   46441: out<=0;
   46442: out<=0;
   46443: out<=1;
   46444: out<=1;
   46445: out<=1;
   46446: out<=1;
   46447: out<=1;
   46448: out<=0;
   46449: out<=0;
   46450: out<=1;
   46451: out<=1;
   46452: out<=0;
   46453: out<=1;
   46454: out<=0;
   46455: out<=1;
   46456: out<=1;
   46457: out<=0;
   46458: out<=0;
   46459: out<=1;
   46460: out<=1;
   46461: out<=1;
   46462: out<=1;
   46463: out<=1;
   46464: out<=1;
   46465: out<=1;
   46466: out<=0;
   46467: out<=0;
   46468: out<=1;
   46469: out<=0;
   46470: out<=1;
   46471: out<=0;
   46472: out<=0;
   46473: out<=1;
   46474: out<=1;
   46475: out<=0;
   46476: out<=0;
   46477: out<=0;
   46478: out<=0;
   46479: out<=0;
   46480: out<=1;
   46481: out<=1;
   46482: out<=0;
   46483: out<=0;
   46484: out<=1;
   46485: out<=0;
   46486: out<=1;
   46487: out<=0;
   46488: out<=0;
   46489: out<=1;
   46490: out<=1;
   46491: out<=0;
   46492: out<=0;
   46493: out<=0;
   46494: out<=0;
   46495: out<=0;
   46496: out<=1;
   46497: out<=1;
   46498: out<=0;
   46499: out<=0;
   46500: out<=1;
   46501: out<=0;
   46502: out<=1;
   46503: out<=0;
   46504: out<=0;
   46505: out<=1;
   46506: out<=1;
   46507: out<=0;
   46508: out<=0;
   46509: out<=0;
   46510: out<=0;
   46511: out<=0;
   46512: out<=1;
   46513: out<=1;
   46514: out<=0;
   46515: out<=0;
   46516: out<=1;
   46517: out<=0;
   46518: out<=1;
   46519: out<=0;
   46520: out<=0;
   46521: out<=1;
   46522: out<=1;
   46523: out<=0;
   46524: out<=0;
   46525: out<=0;
   46526: out<=0;
   46527: out<=0;
   46528: out<=0;
   46529: out<=0;
   46530: out<=1;
   46531: out<=1;
   46532: out<=0;
   46533: out<=1;
   46534: out<=0;
   46535: out<=1;
   46536: out<=1;
   46537: out<=0;
   46538: out<=0;
   46539: out<=1;
   46540: out<=1;
   46541: out<=1;
   46542: out<=1;
   46543: out<=1;
   46544: out<=1;
   46545: out<=1;
   46546: out<=0;
   46547: out<=0;
   46548: out<=1;
   46549: out<=0;
   46550: out<=1;
   46551: out<=0;
   46552: out<=0;
   46553: out<=1;
   46554: out<=1;
   46555: out<=0;
   46556: out<=0;
   46557: out<=0;
   46558: out<=0;
   46559: out<=0;
   46560: out<=1;
   46561: out<=1;
   46562: out<=0;
   46563: out<=0;
   46564: out<=1;
   46565: out<=0;
   46566: out<=1;
   46567: out<=0;
   46568: out<=0;
   46569: out<=1;
   46570: out<=1;
   46571: out<=0;
   46572: out<=0;
   46573: out<=0;
   46574: out<=0;
   46575: out<=0;
   46576: out<=0;
   46577: out<=0;
   46578: out<=1;
   46579: out<=1;
   46580: out<=0;
   46581: out<=1;
   46582: out<=0;
   46583: out<=1;
   46584: out<=1;
   46585: out<=0;
   46586: out<=0;
   46587: out<=1;
   46588: out<=1;
   46589: out<=1;
   46590: out<=1;
   46591: out<=1;
   46592: out<=0;
   46593: out<=0;
   46594: out<=0;
   46595: out<=0;
   46596: out<=0;
   46597: out<=1;
   46598: out<=1;
   46599: out<=0;
   46600: out<=0;
   46601: out<=1;
   46602: out<=0;
   46603: out<=1;
   46604: out<=0;
   46605: out<=0;
   46606: out<=1;
   46607: out<=1;
   46608: out<=1;
   46609: out<=1;
   46610: out<=1;
   46611: out<=1;
   46612: out<=1;
   46613: out<=0;
   46614: out<=0;
   46615: out<=1;
   46616: out<=1;
   46617: out<=0;
   46618: out<=1;
   46619: out<=0;
   46620: out<=1;
   46621: out<=1;
   46622: out<=0;
   46623: out<=0;
   46624: out<=1;
   46625: out<=1;
   46626: out<=1;
   46627: out<=1;
   46628: out<=1;
   46629: out<=0;
   46630: out<=0;
   46631: out<=1;
   46632: out<=1;
   46633: out<=0;
   46634: out<=1;
   46635: out<=0;
   46636: out<=1;
   46637: out<=1;
   46638: out<=0;
   46639: out<=0;
   46640: out<=0;
   46641: out<=0;
   46642: out<=0;
   46643: out<=0;
   46644: out<=0;
   46645: out<=1;
   46646: out<=1;
   46647: out<=0;
   46648: out<=0;
   46649: out<=1;
   46650: out<=0;
   46651: out<=1;
   46652: out<=0;
   46653: out<=0;
   46654: out<=1;
   46655: out<=1;
   46656: out<=1;
   46657: out<=1;
   46658: out<=1;
   46659: out<=1;
   46660: out<=1;
   46661: out<=0;
   46662: out<=0;
   46663: out<=1;
   46664: out<=1;
   46665: out<=0;
   46666: out<=1;
   46667: out<=0;
   46668: out<=1;
   46669: out<=1;
   46670: out<=0;
   46671: out<=0;
   46672: out<=1;
   46673: out<=1;
   46674: out<=1;
   46675: out<=1;
   46676: out<=1;
   46677: out<=0;
   46678: out<=0;
   46679: out<=1;
   46680: out<=1;
   46681: out<=0;
   46682: out<=1;
   46683: out<=0;
   46684: out<=1;
   46685: out<=1;
   46686: out<=0;
   46687: out<=0;
   46688: out<=1;
   46689: out<=1;
   46690: out<=1;
   46691: out<=1;
   46692: out<=1;
   46693: out<=0;
   46694: out<=0;
   46695: out<=1;
   46696: out<=1;
   46697: out<=0;
   46698: out<=1;
   46699: out<=0;
   46700: out<=1;
   46701: out<=1;
   46702: out<=0;
   46703: out<=0;
   46704: out<=1;
   46705: out<=1;
   46706: out<=1;
   46707: out<=1;
   46708: out<=1;
   46709: out<=0;
   46710: out<=0;
   46711: out<=1;
   46712: out<=1;
   46713: out<=0;
   46714: out<=1;
   46715: out<=0;
   46716: out<=1;
   46717: out<=1;
   46718: out<=0;
   46719: out<=0;
   46720: out<=1;
   46721: out<=1;
   46722: out<=1;
   46723: out<=1;
   46724: out<=1;
   46725: out<=0;
   46726: out<=0;
   46727: out<=1;
   46728: out<=1;
   46729: out<=0;
   46730: out<=1;
   46731: out<=0;
   46732: out<=1;
   46733: out<=1;
   46734: out<=0;
   46735: out<=0;
   46736: out<=1;
   46737: out<=1;
   46738: out<=1;
   46739: out<=1;
   46740: out<=1;
   46741: out<=0;
   46742: out<=0;
   46743: out<=1;
   46744: out<=1;
   46745: out<=0;
   46746: out<=1;
   46747: out<=0;
   46748: out<=1;
   46749: out<=1;
   46750: out<=0;
   46751: out<=0;
   46752: out<=0;
   46753: out<=0;
   46754: out<=0;
   46755: out<=0;
   46756: out<=0;
   46757: out<=1;
   46758: out<=1;
   46759: out<=0;
   46760: out<=0;
   46761: out<=1;
   46762: out<=0;
   46763: out<=1;
   46764: out<=0;
   46765: out<=0;
   46766: out<=1;
   46767: out<=1;
   46768: out<=0;
   46769: out<=0;
   46770: out<=0;
   46771: out<=0;
   46772: out<=0;
   46773: out<=1;
   46774: out<=1;
   46775: out<=0;
   46776: out<=0;
   46777: out<=1;
   46778: out<=0;
   46779: out<=1;
   46780: out<=0;
   46781: out<=0;
   46782: out<=1;
   46783: out<=1;
   46784: out<=0;
   46785: out<=0;
   46786: out<=0;
   46787: out<=0;
   46788: out<=0;
   46789: out<=1;
   46790: out<=1;
   46791: out<=0;
   46792: out<=0;
   46793: out<=1;
   46794: out<=0;
   46795: out<=1;
   46796: out<=0;
   46797: out<=0;
   46798: out<=1;
   46799: out<=1;
   46800: out<=1;
   46801: out<=1;
   46802: out<=1;
   46803: out<=1;
   46804: out<=1;
   46805: out<=0;
   46806: out<=0;
   46807: out<=1;
   46808: out<=1;
   46809: out<=0;
   46810: out<=1;
   46811: out<=0;
   46812: out<=1;
   46813: out<=1;
   46814: out<=0;
   46815: out<=0;
   46816: out<=0;
   46817: out<=0;
   46818: out<=0;
   46819: out<=0;
   46820: out<=0;
   46821: out<=1;
   46822: out<=1;
   46823: out<=0;
   46824: out<=0;
   46825: out<=1;
   46826: out<=0;
   46827: out<=1;
   46828: out<=0;
   46829: out<=0;
   46830: out<=1;
   46831: out<=1;
   46832: out<=1;
   46833: out<=1;
   46834: out<=1;
   46835: out<=1;
   46836: out<=1;
   46837: out<=0;
   46838: out<=0;
   46839: out<=1;
   46840: out<=1;
   46841: out<=0;
   46842: out<=1;
   46843: out<=0;
   46844: out<=1;
   46845: out<=1;
   46846: out<=0;
   46847: out<=0;
   46848: out<=1;
   46849: out<=0;
   46850: out<=0;
   46851: out<=1;
   46852: out<=0;
   46853: out<=0;
   46854: out<=0;
   46855: out<=0;
   46856: out<=0;
   46857: out<=0;
   46858: out<=1;
   46859: out<=1;
   46860: out<=1;
   46861: out<=0;
   46862: out<=1;
   46863: out<=0;
   46864: out<=1;
   46865: out<=0;
   46866: out<=0;
   46867: out<=1;
   46868: out<=0;
   46869: out<=0;
   46870: out<=0;
   46871: out<=0;
   46872: out<=0;
   46873: out<=0;
   46874: out<=1;
   46875: out<=1;
   46876: out<=1;
   46877: out<=0;
   46878: out<=1;
   46879: out<=0;
   46880: out<=1;
   46881: out<=0;
   46882: out<=0;
   46883: out<=1;
   46884: out<=0;
   46885: out<=0;
   46886: out<=0;
   46887: out<=0;
   46888: out<=0;
   46889: out<=0;
   46890: out<=1;
   46891: out<=1;
   46892: out<=1;
   46893: out<=0;
   46894: out<=1;
   46895: out<=0;
   46896: out<=1;
   46897: out<=0;
   46898: out<=0;
   46899: out<=1;
   46900: out<=0;
   46901: out<=0;
   46902: out<=0;
   46903: out<=0;
   46904: out<=0;
   46905: out<=0;
   46906: out<=1;
   46907: out<=1;
   46908: out<=1;
   46909: out<=0;
   46910: out<=1;
   46911: out<=0;
   46912: out<=0;
   46913: out<=1;
   46914: out<=1;
   46915: out<=0;
   46916: out<=1;
   46917: out<=1;
   46918: out<=1;
   46919: out<=1;
   46920: out<=1;
   46921: out<=1;
   46922: out<=0;
   46923: out<=0;
   46924: out<=0;
   46925: out<=1;
   46926: out<=0;
   46927: out<=1;
   46928: out<=1;
   46929: out<=0;
   46930: out<=0;
   46931: out<=1;
   46932: out<=0;
   46933: out<=0;
   46934: out<=0;
   46935: out<=0;
   46936: out<=0;
   46937: out<=0;
   46938: out<=1;
   46939: out<=1;
   46940: out<=1;
   46941: out<=0;
   46942: out<=1;
   46943: out<=0;
   46944: out<=1;
   46945: out<=0;
   46946: out<=0;
   46947: out<=1;
   46948: out<=0;
   46949: out<=0;
   46950: out<=0;
   46951: out<=0;
   46952: out<=0;
   46953: out<=0;
   46954: out<=1;
   46955: out<=1;
   46956: out<=1;
   46957: out<=0;
   46958: out<=1;
   46959: out<=0;
   46960: out<=0;
   46961: out<=1;
   46962: out<=1;
   46963: out<=0;
   46964: out<=1;
   46965: out<=1;
   46966: out<=1;
   46967: out<=1;
   46968: out<=1;
   46969: out<=1;
   46970: out<=0;
   46971: out<=0;
   46972: out<=0;
   46973: out<=1;
   46974: out<=0;
   46975: out<=1;
   46976: out<=0;
   46977: out<=1;
   46978: out<=1;
   46979: out<=0;
   46980: out<=1;
   46981: out<=1;
   46982: out<=1;
   46983: out<=1;
   46984: out<=1;
   46985: out<=1;
   46986: out<=0;
   46987: out<=0;
   46988: out<=0;
   46989: out<=1;
   46990: out<=0;
   46991: out<=1;
   46992: out<=1;
   46993: out<=0;
   46994: out<=0;
   46995: out<=1;
   46996: out<=0;
   46997: out<=0;
   46998: out<=0;
   46999: out<=0;
   47000: out<=0;
   47001: out<=0;
   47002: out<=1;
   47003: out<=1;
   47004: out<=1;
   47005: out<=0;
   47006: out<=1;
   47007: out<=0;
   47008: out<=0;
   47009: out<=1;
   47010: out<=1;
   47011: out<=0;
   47012: out<=1;
   47013: out<=1;
   47014: out<=1;
   47015: out<=1;
   47016: out<=1;
   47017: out<=1;
   47018: out<=0;
   47019: out<=0;
   47020: out<=0;
   47021: out<=1;
   47022: out<=0;
   47023: out<=1;
   47024: out<=1;
   47025: out<=0;
   47026: out<=0;
   47027: out<=1;
   47028: out<=0;
   47029: out<=0;
   47030: out<=0;
   47031: out<=0;
   47032: out<=0;
   47033: out<=0;
   47034: out<=1;
   47035: out<=1;
   47036: out<=1;
   47037: out<=0;
   47038: out<=1;
   47039: out<=0;
   47040: out<=1;
   47041: out<=0;
   47042: out<=0;
   47043: out<=1;
   47044: out<=0;
   47045: out<=0;
   47046: out<=0;
   47047: out<=0;
   47048: out<=0;
   47049: out<=0;
   47050: out<=1;
   47051: out<=1;
   47052: out<=1;
   47053: out<=0;
   47054: out<=1;
   47055: out<=0;
   47056: out<=1;
   47057: out<=0;
   47058: out<=0;
   47059: out<=1;
   47060: out<=0;
   47061: out<=0;
   47062: out<=0;
   47063: out<=0;
   47064: out<=0;
   47065: out<=0;
   47066: out<=1;
   47067: out<=1;
   47068: out<=1;
   47069: out<=0;
   47070: out<=1;
   47071: out<=0;
   47072: out<=0;
   47073: out<=1;
   47074: out<=1;
   47075: out<=0;
   47076: out<=1;
   47077: out<=1;
   47078: out<=1;
   47079: out<=1;
   47080: out<=1;
   47081: out<=1;
   47082: out<=0;
   47083: out<=0;
   47084: out<=0;
   47085: out<=1;
   47086: out<=0;
   47087: out<=1;
   47088: out<=0;
   47089: out<=1;
   47090: out<=1;
   47091: out<=0;
   47092: out<=1;
   47093: out<=1;
   47094: out<=1;
   47095: out<=1;
   47096: out<=1;
   47097: out<=1;
   47098: out<=0;
   47099: out<=0;
   47100: out<=0;
   47101: out<=1;
   47102: out<=0;
   47103: out<=1;
   47104: out<=1;
   47105: out<=0;
   47106: out<=0;
   47107: out<=1;
   47108: out<=0;
   47109: out<=0;
   47110: out<=0;
   47111: out<=0;
   47112: out<=1;
   47113: out<=1;
   47114: out<=0;
   47115: out<=0;
   47116: out<=0;
   47117: out<=1;
   47118: out<=0;
   47119: out<=1;
   47120: out<=1;
   47121: out<=0;
   47122: out<=0;
   47123: out<=1;
   47124: out<=0;
   47125: out<=0;
   47126: out<=0;
   47127: out<=0;
   47128: out<=1;
   47129: out<=1;
   47130: out<=0;
   47131: out<=0;
   47132: out<=0;
   47133: out<=1;
   47134: out<=0;
   47135: out<=1;
   47136: out<=0;
   47137: out<=1;
   47138: out<=1;
   47139: out<=0;
   47140: out<=1;
   47141: out<=1;
   47142: out<=1;
   47143: out<=1;
   47144: out<=0;
   47145: out<=0;
   47146: out<=1;
   47147: out<=1;
   47148: out<=1;
   47149: out<=0;
   47150: out<=1;
   47151: out<=0;
   47152: out<=0;
   47153: out<=1;
   47154: out<=1;
   47155: out<=0;
   47156: out<=1;
   47157: out<=1;
   47158: out<=1;
   47159: out<=1;
   47160: out<=0;
   47161: out<=0;
   47162: out<=1;
   47163: out<=1;
   47164: out<=1;
   47165: out<=0;
   47166: out<=1;
   47167: out<=0;
   47168: out<=0;
   47169: out<=1;
   47170: out<=1;
   47171: out<=0;
   47172: out<=1;
   47173: out<=1;
   47174: out<=1;
   47175: out<=1;
   47176: out<=0;
   47177: out<=0;
   47178: out<=1;
   47179: out<=1;
   47180: out<=1;
   47181: out<=0;
   47182: out<=1;
   47183: out<=0;
   47184: out<=1;
   47185: out<=0;
   47186: out<=0;
   47187: out<=1;
   47188: out<=0;
   47189: out<=0;
   47190: out<=0;
   47191: out<=0;
   47192: out<=1;
   47193: out<=1;
   47194: out<=0;
   47195: out<=0;
   47196: out<=0;
   47197: out<=1;
   47198: out<=0;
   47199: out<=1;
   47200: out<=0;
   47201: out<=1;
   47202: out<=1;
   47203: out<=0;
   47204: out<=1;
   47205: out<=1;
   47206: out<=1;
   47207: out<=1;
   47208: out<=0;
   47209: out<=0;
   47210: out<=1;
   47211: out<=1;
   47212: out<=1;
   47213: out<=0;
   47214: out<=1;
   47215: out<=0;
   47216: out<=1;
   47217: out<=0;
   47218: out<=0;
   47219: out<=1;
   47220: out<=0;
   47221: out<=0;
   47222: out<=0;
   47223: out<=0;
   47224: out<=1;
   47225: out<=1;
   47226: out<=0;
   47227: out<=0;
   47228: out<=0;
   47229: out<=1;
   47230: out<=0;
   47231: out<=1;
   47232: out<=0;
   47233: out<=1;
   47234: out<=1;
   47235: out<=0;
   47236: out<=1;
   47237: out<=1;
   47238: out<=1;
   47239: out<=1;
   47240: out<=0;
   47241: out<=0;
   47242: out<=1;
   47243: out<=1;
   47244: out<=1;
   47245: out<=0;
   47246: out<=1;
   47247: out<=0;
   47248: out<=1;
   47249: out<=0;
   47250: out<=0;
   47251: out<=1;
   47252: out<=0;
   47253: out<=0;
   47254: out<=0;
   47255: out<=0;
   47256: out<=1;
   47257: out<=1;
   47258: out<=0;
   47259: out<=0;
   47260: out<=0;
   47261: out<=1;
   47262: out<=0;
   47263: out<=1;
   47264: out<=1;
   47265: out<=0;
   47266: out<=0;
   47267: out<=1;
   47268: out<=0;
   47269: out<=0;
   47270: out<=0;
   47271: out<=0;
   47272: out<=1;
   47273: out<=1;
   47274: out<=0;
   47275: out<=0;
   47276: out<=0;
   47277: out<=1;
   47278: out<=0;
   47279: out<=1;
   47280: out<=0;
   47281: out<=1;
   47282: out<=1;
   47283: out<=0;
   47284: out<=1;
   47285: out<=1;
   47286: out<=1;
   47287: out<=1;
   47288: out<=0;
   47289: out<=0;
   47290: out<=1;
   47291: out<=1;
   47292: out<=1;
   47293: out<=0;
   47294: out<=1;
   47295: out<=0;
   47296: out<=1;
   47297: out<=0;
   47298: out<=0;
   47299: out<=1;
   47300: out<=0;
   47301: out<=0;
   47302: out<=0;
   47303: out<=0;
   47304: out<=1;
   47305: out<=1;
   47306: out<=0;
   47307: out<=0;
   47308: out<=0;
   47309: out<=1;
   47310: out<=0;
   47311: out<=1;
   47312: out<=1;
   47313: out<=0;
   47314: out<=0;
   47315: out<=1;
   47316: out<=0;
   47317: out<=0;
   47318: out<=0;
   47319: out<=0;
   47320: out<=1;
   47321: out<=1;
   47322: out<=0;
   47323: out<=0;
   47324: out<=0;
   47325: out<=1;
   47326: out<=0;
   47327: out<=1;
   47328: out<=1;
   47329: out<=0;
   47330: out<=0;
   47331: out<=1;
   47332: out<=0;
   47333: out<=0;
   47334: out<=0;
   47335: out<=0;
   47336: out<=1;
   47337: out<=1;
   47338: out<=0;
   47339: out<=0;
   47340: out<=0;
   47341: out<=1;
   47342: out<=0;
   47343: out<=1;
   47344: out<=1;
   47345: out<=0;
   47346: out<=0;
   47347: out<=1;
   47348: out<=0;
   47349: out<=0;
   47350: out<=0;
   47351: out<=0;
   47352: out<=1;
   47353: out<=1;
   47354: out<=0;
   47355: out<=0;
   47356: out<=0;
   47357: out<=1;
   47358: out<=0;
   47359: out<=1;
   47360: out<=0;
   47361: out<=0;
   47362: out<=0;
   47363: out<=0;
   47364: out<=0;
   47365: out<=1;
   47366: out<=1;
   47367: out<=0;
   47368: out<=1;
   47369: out<=0;
   47370: out<=1;
   47371: out<=0;
   47372: out<=1;
   47373: out<=1;
   47374: out<=0;
   47375: out<=0;
   47376: out<=1;
   47377: out<=1;
   47378: out<=1;
   47379: out<=1;
   47380: out<=1;
   47381: out<=0;
   47382: out<=0;
   47383: out<=1;
   47384: out<=0;
   47385: out<=1;
   47386: out<=0;
   47387: out<=1;
   47388: out<=0;
   47389: out<=0;
   47390: out<=1;
   47391: out<=1;
   47392: out<=0;
   47393: out<=0;
   47394: out<=0;
   47395: out<=0;
   47396: out<=0;
   47397: out<=1;
   47398: out<=1;
   47399: out<=0;
   47400: out<=1;
   47401: out<=0;
   47402: out<=1;
   47403: out<=0;
   47404: out<=1;
   47405: out<=1;
   47406: out<=0;
   47407: out<=0;
   47408: out<=1;
   47409: out<=1;
   47410: out<=1;
   47411: out<=1;
   47412: out<=1;
   47413: out<=0;
   47414: out<=0;
   47415: out<=1;
   47416: out<=0;
   47417: out<=1;
   47418: out<=0;
   47419: out<=1;
   47420: out<=0;
   47421: out<=0;
   47422: out<=1;
   47423: out<=1;
   47424: out<=1;
   47425: out<=1;
   47426: out<=1;
   47427: out<=1;
   47428: out<=1;
   47429: out<=0;
   47430: out<=0;
   47431: out<=1;
   47432: out<=0;
   47433: out<=1;
   47434: out<=0;
   47435: out<=1;
   47436: out<=0;
   47437: out<=0;
   47438: out<=1;
   47439: out<=1;
   47440: out<=1;
   47441: out<=1;
   47442: out<=1;
   47443: out<=1;
   47444: out<=1;
   47445: out<=0;
   47446: out<=0;
   47447: out<=1;
   47448: out<=0;
   47449: out<=1;
   47450: out<=0;
   47451: out<=1;
   47452: out<=0;
   47453: out<=0;
   47454: out<=1;
   47455: out<=1;
   47456: out<=0;
   47457: out<=0;
   47458: out<=0;
   47459: out<=0;
   47460: out<=0;
   47461: out<=1;
   47462: out<=1;
   47463: out<=0;
   47464: out<=1;
   47465: out<=0;
   47466: out<=1;
   47467: out<=0;
   47468: out<=1;
   47469: out<=1;
   47470: out<=0;
   47471: out<=0;
   47472: out<=0;
   47473: out<=0;
   47474: out<=0;
   47475: out<=0;
   47476: out<=0;
   47477: out<=1;
   47478: out<=1;
   47479: out<=0;
   47480: out<=1;
   47481: out<=0;
   47482: out<=1;
   47483: out<=0;
   47484: out<=1;
   47485: out<=1;
   47486: out<=0;
   47487: out<=0;
   47488: out<=1;
   47489: out<=1;
   47490: out<=1;
   47491: out<=1;
   47492: out<=1;
   47493: out<=0;
   47494: out<=0;
   47495: out<=1;
   47496: out<=0;
   47497: out<=1;
   47498: out<=0;
   47499: out<=1;
   47500: out<=0;
   47501: out<=0;
   47502: out<=1;
   47503: out<=1;
   47504: out<=1;
   47505: out<=1;
   47506: out<=1;
   47507: out<=1;
   47508: out<=1;
   47509: out<=0;
   47510: out<=0;
   47511: out<=1;
   47512: out<=0;
   47513: out<=1;
   47514: out<=0;
   47515: out<=1;
   47516: out<=0;
   47517: out<=0;
   47518: out<=1;
   47519: out<=1;
   47520: out<=1;
   47521: out<=1;
   47522: out<=1;
   47523: out<=1;
   47524: out<=1;
   47525: out<=0;
   47526: out<=0;
   47527: out<=1;
   47528: out<=0;
   47529: out<=1;
   47530: out<=0;
   47531: out<=1;
   47532: out<=0;
   47533: out<=0;
   47534: out<=1;
   47535: out<=1;
   47536: out<=1;
   47537: out<=1;
   47538: out<=1;
   47539: out<=1;
   47540: out<=1;
   47541: out<=0;
   47542: out<=0;
   47543: out<=1;
   47544: out<=0;
   47545: out<=1;
   47546: out<=0;
   47547: out<=1;
   47548: out<=0;
   47549: out<=0;
   47550: out<=1;
   47551: out<=1;
   47552: out<=0;
   47553: out<=0;
   47554: out<=0;
   47555: out<=0;
   47556: out<=0;
   47557: out<=1;
   47558: out<=1;
   47559: out<=0;
   47560: out<=1;
   47561: out<=0;
   47562: out<=1;
   47563: out<=0;
   47564: out<=1;
   47565: out<=1;
   47566: out<=0;
   47567: out<=0;
   47568: out<=1;
   47569: out<=1;
   47570: out<=1;
   47571: out<=1;
   47572: out<=1;
   47573: out<=0;
   47574: out<=0;
   47575: out<=1;
   47576: out<=0;
   47577: out<=1;
   47578: out<=0;
   47579: out<=1;
   47580: out<=0;
   47581: out<=0;
   47582: out<=1;
   47583: out<=1;
   47584: out<=1;
   47585: out<=1;
   47586: out<=1;
   47587: out<=1;
   47588: out<=1;
   47589: out<=0;
   47590: out<=0;
   47591: out<=1;
   47592: out<=0;
   47593: out<=1;
   47594: out<=0;
   47595: out<=1;
   47596: out<=0;
   47597: out<=0;
   47598: out<=1;
   47599: out<=1;
   47600: out<=0;
   47601: out<=0;
   47602: out<=0;
   47603: out<=0;
   47604: out<=0;
   47605: out<=1;
   47606: out<=1;
   47607: out<=0;
   47608: out<=1;
   47609: out<=0;
   47610: out<=1;
   47611: out<=0;
   47612: out<=1;
   47613: out<=1;
   47614: out<=0;
   47615: out<=0;
   47616: out<=1;
   47617: out<=1;
   47618: out<=0;
   47619: out<=0;
   47620: out<=1;
   47621: out<=0;
   47622: out<=1;
   47623: out<=0;
   47624: out<=1;
   47625: out<=0;
   47626: out<=0;
   47627: out<=1;
   47628: out<=1;
   47629: out<=1;
   47630: out<=1;
   47631: out<=1;
   47632: out<=0;
   47633: out<=0;
   47634: out<=1;
   47635: out<=1;
   47636: out<=0;
   47637: out<=1;
   47638: out<=0;
   47639: out<=1;
   47640: out<=0;
   47641: out<=1;
   47642: out<=1;
   47643: out<=0;
   47644: out<=0;
   47645: out<=0;
   47646: out<=0;
   47647: out<=0;
   47648: out<=0;
   47649: out<=0;
   47650: out<=1;
   47651: out<=1;
   47652: out<=0;
   47653: out<=1;
   47654: out<=0;
   47655: out<=1;
   47656: out<=0;
   47657: out<=1;
   47658: out<=1;
   47659: out<=0;
   47660: out<=0;
   47661: out<=0;
   47662: out<=0;
   47663: out<=0;
   47664: out<=1;
   47665: out<=1;
   47666: out<=0;
   47667: out<=0;
   47668: out<=1;
   47669: out<=0;
   47670: out<=1;
   47671: out<=0;
   47672: out<=1;
   47673: out<=0;
   47674: out<=0;
   47675: out<=1;
   47676: out<=1;
   47677: out<=1;
   47678: out<=1;
   47679: out<=1;
   47680: out<=0;
   47681: out<=0;
   47682: out<=1;
   47683: out<=1;
   47684: out<=0;
   47685: out<=1;
   47686: out<=0;
   47687: out<=1;
   47688: out<=0;
   47689: out<=1;
   47690: out<=1;
   47691: out<=0;
   47692: out<=0;
   47693: out<=0;
   47694: out<=0;
   47695: out<=0;
   47696: out<=0;
   47697: out<=0;
   47698: out<=1;
   47699: out<=1;
   47700: out<=0;
   47701: out<=1;
   47702: out<=0;
   47703: out<=1;
   47704: out<=0;
   47705: out<=1;
   47706: out<=1;
   47707: out<=0;
   47708: out<=0;
   47709: out<=0;
   47710: out<=0;
   47711: out<=0;
   47712: out<=0;
   47713: out<=0;
   47714: out<=1;
   47715: out<=1;
   47716: out<=0;
   47717: out<=1;
   47718: out<=0;
   47719: out<=1;
   47720: out<=0;
   47721: out<=1;
   47722: out<=1;
   47723: out<=0;
   47724: out<=0;
   47725: out<=0;
   47726: out<=0;
   47727: out<=0;
   47728: out<=0;
   47729: out<=0;
   47730: out<=1;
   47731: out<=1;
   47732: out<=0;
   47733: out<=1;
   47734: out<=0;
   47735: out<=1;
   47736: out<=0;
   47737: out<=1;
   47738: out<=1;
   47739: out<=0;
   47740: out<=0;
   47741: out<=0;
   47742: out<=0;
   47743: out<=0;
   47744: out<=0;
   47745: out<=0;
   47746: out<=1;
   47747: out<=1;
   47748: out<=0;
   47749: out<=1;
   47750: out<=0;
   47751: out<=1;
   47752: out<=0;
   47753: out<=1;
   47754: out<=1;
   47755: out<=0;
   47756: out<=0;
   47757: out<=0;
   47758: out<=0;
   47759: out<=0;
   47760: out<=0;
   47761: out<=0;
   47762: out<=1;
   47763: out<=1;
   47764: out<=0;
   47765: out<=1;
   47766: out<=0;
   47767: out<=1;
   47768: out<=0;
   47769: out<=1;
   47770: out<=1;
   47771: out<=0;
   47772: out<=0;
   47773: out<=0;
   47774: out<=0;
   47775: out<=0;
   47776: out<=1;
   47777: out<=1;
   47778: out<=0;
   47779: out<=0;
   47780: out<=1;
   47781: out<=0;
   47782: out<=1;
   47783: out<=0;
   47784: out<=1;
   47785: out<=0;
   47786: out<=0;
   47787: out<=1;
   47788: out<=1;
   47789: out<=1;
   47790: out<=1;
   47791: out<=1;
   47792: out<=1;
   47793: out<=1;
   47794: out<=0;
   47795: out<=0;
   47796: out<=1;
   47797: out<=0;
   47798: out<=1;
   47799: out<=0;
   47800: out<=1;
   47801: out<=0;
   47802: out<=0;
   47803: out<=1;
   47804: out<=1;
   47805: out<=1;
   47806: out<=1;
   47807: out<=1;
   47808: out<=1;
   47809: out<=1;
   47810: out<=0;
   47811: out<=0;
   47812: out<=1;
   47813: out<=0;
   47814: out<=1;
   47815: out<=0;
   47816: out<=1;
   47817: out<=0;
   47818: out<=0;
   47819: out<=1;
   47820: out<=1;
   47821: out<=1;
   47822: out<=1;
   47823: out<=1;
   47824: out<=0;
   47825: out<=0;
   47826: out<=1;
   47827: out<=1;
   47828: out<=0;
   47829: out<=1;
   47830: out<=0;
   47831: out<=1;
   47832: out<=0;
   47833: out<=1;
   47834: out<=1;
   47835: out<=0;
   47836: out<=0;
   47837: out<=0;
   47838: out<=0;
   47839: out<=0;
   47840: out<=1;
   47841: out<=1;
   47842: out<=0;
   47843: out<=0;
   47844: out<=1;
   47845: out<=0;
   47846: out<=1;
   47847: out<=0;
   47848: out<=1;
   47849: out<=0;
   47850: out<=0;
   47851: out<=1;
   47852: out<=1;
   47853: out<=1;
   47854: out<=1;
   47855: out<=1;
   47856: out<=0;
   47857: out<=0;
   47858: out<=1;
   47859: out<=1;
   47860: out<=0;
   47861: out<=1;
   47862: out<=0;
   47863: out<=1;
   47864: out<=0;
   47865: out<=1;
   47866: out<=1;
   47867: out<=0;
   47868: out<=0;
   47869: out<=0;
   47870: out<=0;
   47871: out<=0;
   47872: out<=0;
   47873: out<=1;
   47874: out<=0;
   47875: out<=1;
   47876: out<=1;
   47877: out<=1;
   47878: out<=0;
   47879: out<=0;
   47880: out<=1;
   47881: out<=1;
   47882: out<=1;
   47883: out<=1;
   47884: out<=0;
   47885: out<=1;
   47886: out<=1;
   47887: out<=0;
   47888: out<=0;
   47889: out<=1;
   47890: out<=0;
   47891: out<=1;
   47892: out<=1;
   47893: out<=1;
   47894: out<=0;
   47895: out<=0;
   47896: out<=1;
   47897: out<=1;
   47898: out<=1;
   47899: out<=1;
   47900: out<=0;
   47901: out<=1;
   47902: out<=1;
   47903: out<=0;
   47904: out<=0;
   47905: out<=1;
   47906: out<=0;
   47907: out<=1;
   47908: out<=1;
   47909: out<=1;
   47910: out<=0;
   47911: out<=0;
   47912: out<=1;
   47913: out<=1;
   47914: out<=1;
   47915: out<=1;
   47916: out<=0;
   47917: out<=1;
   47918: out<=1;
   47919: out<=0;
   47920: out<=0;
   47921: out<=1;
   47922: out<=0;
   47923: out<=1;
   47924: out<=1;
   47925: out<=1;
   47926: out<=0;
   47927: out<=0;
   47928: out<=1;
   47929: out<=1;
   47930: out<=1;
   47931: out<=1;
   47932: out<=0;
   47933: out<=1;
   47934: out<=1;
   47935: out<=0;
   47936: out<=1;
   47937: out<=0;
   47938: out<=1;
   47939: out<=0;
   47940: out<=0;
   47941: out<=0;
   47942: out<=1;
   47943: out<=1;
   47944: out<=0;
   47945: out<=0;
   47946: out<=0;
   47947: out<=0;
   47948: out<=1;
   47949: out<=0;
   47950: out<=0;
   47951: out<=1;
   47952: out<=0;
   47953: out<=1;
   47954: out<=0;
   47955: out<=1;
   47956: out<=1;
   47957: out<=1;
   47958: out<=0;
   47959: out<=0;
   47960: out<=1;
   47961: out<=1;
   47962: out<=1;
   47963: out<=1;
   47964: out<=0;
   47965: out<=1;
   47966: out<=1;
   47967: out<=0;
   47968: out<=0;
   47969: out<=1;
   47970: out<=0;
   47971: out<=1;
   47972: out<=1;
   47973: out<=1;
   47974: out<=0;
   47975: out<=0;
   47976: out<=1;
   47977: out<=1;
   47978: out<=1;
   47979: out<=1;
   47980: out<=0;
   47981: out<=1;
   47982: out<=1;
   47983: out<=0;
   47984: out<=1;
   47985: out<=0;
   47986: out<=1;
   47987: out<=0;
   47988: out<=0;
   47989: out<=0;
   47990: out<=1;
   47991: out<=1;
   47992: out<=0;
   47993: out<=0;
   47994: out<=0;
   47995: out<=0;
   47996: out<=1;
   47997: out<=0;
   47998: out<=0;
   47999: out<=1;
   48000: out<=1;
   48001: out<=0;
   48002: out<=1;
   48003: out<=0;
   48004: out<=0;
   48005: out<=0;
   48006: out<=1;
   48007: out<=1;
   48008: out<=0;
   48009: out<=0;
   48010: out<=0;
   48011: out<=0;
   48012: out<=1;
   48013: out<=0;
   48014: out<=0;
   48015: out<=1;
   48016: out<=0;
   48017: out<=1;
   48018: out<=0;
   48019: out<=1;
   48020: out<=1;
   48021: out<=1;
   48022: out<=0;
   48023: out<=0;
   48024: out<=1;
   48025: out<=1;
   48026: out<=1;
   48027: out<=1;
   48028: out<=0;
   48029: out<=1;
   48030: out<=1;
   48031: out<=0;
   48032: out<=1;
   48033: out<=0;
   48034: out<=1;
   48035: out<=0;
   48036: out<=0;
   48037: out<=0;
   48038: out<=1;
   48039: out<=1;
   48040: out<=0;
   48041: out<=0;
   48042: out<=0;
   48043: out<=0;
   48044: out<=1;
   48045: out<=0;
   48046: out<=0;
   48047: out<=1;
   48048: out<=0;
   48049: out<=1;
   48050: out<=0;
   48051: out<=1;
   48052: out<=1;
   48053: out<=1;
   48054: out<=0;
   48055: out<=0;
   48056: out<=1;
   48057: out<=1;
   48058: out<=1;
   48059: out<=1;
   48060: out<=0;
   48061: out<=1;
   48062: out<=1;
   48063: out<=0;
   48064: out<=0;
   48065: out<=1;
   48066: out<=0;
   48067: out<=1;
   48068: out<=1;
   48069: out<=1;
   48070: out<=0;
   48071: out<=0;
   48072: out<=1;
   48073: out<=1;
   48074: out<=1;
   48075: out<=1;
   48076: out<=0;
   48077: out<=1;
   48078: out<=1;
   48079: out<=0;
   48080: out<=0;
   48081: out<=1;
   48082: out<=0;
   48083: out<=1;
   48084: out<=1;
   48085: out<=1;
   48086: out<=0;
   48087: out<=0;
   48088: out<=1;
   48089: out<=1;
   48090: out<=1;
   48091: out<=1;
   48092: out<=0;
   48093: out<=1;
   48094: out<=1;
   48095: out<=0;
   48096: out<=1;
   48097: out<=0;
   48098: out<=1;
   48099: out<=0;
   48100: out<=0;
   48101: out<=0;
   48102: out<=1;
   48103: out<=1;
   48104: out<=0;
   48105: out<=0;
   48106: out<=0;
   48107: out<=0;
   48108: out<=1;
   48109: out<=0;
   48110: out<=0;
   48111: out<=1;
   48112: out<=1;
   48113: out<=0;
   48114: out<=1;
   48115: out<=0;
   48116: out<=0;
   48117: out<=0;
   48118: out<=1;
   48119: out<=1;
   48120: out<=0;
   48121: out<=0;
   48122: out<=0;
   48123: out<=0;
   48124: out<=1;
   48125: out<=0;
   48126: out<=0;
   48127: out<=1;
   48128: out<=1;
   48129: out<=1;
   48130: out<=1;
   48131: out<=1;
   48132: out<=0;
   48133: out<=1;
   48134: out<=1;
   48135: out<=0;
   48136: out<=1;
   48137: out<=0;
   48138: out<=1;
   48139: out<=0;
   48140: out<=0;
   48141: out<=0;
   48142: out<=1;
   48143: out<=1;
   48144: out<=1;
   48145: out<=1;
   48146: out<=1;
   48147: out<=1;
   48148: out<=0;
   48149: out<=1;
   48150: out<=1;
   48151: out<=0;
   48152: out<=1;
   48153: out<=0;
   48154: out<=1;
   48155: out<=0;
   48156: out<=0;
   48157: out<=0;
   48158: out<=1;
   48159: out<=1;
   48160: out<=0;
   48161: out<=0;
   48162: out<=0;
   48163: out<=0;
   48164: out<=1;
   48165: out<=0;
   48166: out<=0;
   48167: out<=1;
   48168: out<=0;
   48169: out<=1;
   48170: out<=0;
   48171: out<=1;
   48172: out<=1;
   48173: out<=1;
   48174: out<=0;
   48175: out<=0;
   48176: out<=0;
   48177: out<=0;
   48178: out<=0;
   48179: out<=0;
   48180: out<=1;
   48181: out<=0;
   48182: out<=0;
   48183: out<=1;
   48184: out<=0;
   48185: out<=1;
   48186: out<=0;
   48187: out<=1;
   48188: out<=1;
   48189: out<=1;
   48190: out<=0;
   48191: out<=0;
   48192: out<=0;
   48193: out<=0;
   48194: out<=0;
   48195: out<=0;
   48196: out<=1;
   48197: out<=0;
   48198: out<=0;
   48199: out<=1;
   48200: out<=0;
   48201: out<=1;
   48202: out<=0;
   48203: out<=1;
   48204: out<=1;
   48205: out<=1;
   48206: out<=0;
   48207: out<=0;
   48208: out<=1;
   48209: out<=1;
   48210: out<=1;
   48211: out<=1;
   48212: out<=0;
   48213: out<=1;
   48214: out<=1;
   48215: out<=0;
   48216: out<=1;
   48217: out<=0;
   48218: out<=1;
   48219: out<=0;
   48220: out<=0;
   48221: out<=0;
   48222: out<=1;
   48223: out<=1;
   48224: out<=0;
   48225: out<=0;
   48226: out<=0;
   48227: out<=0;
   48228: out<=1;
   48229: out<=0;
   48230: out<=0;
   48231: out<=1;
   48232: out<=0;
   48233: out<=1;
   48234: out<=0;
   48235: out<=1;
   48236: out<=1;
   48237: out<=1;
   48238: out<=0;
   48239: out<=0;
   48240: out<=1;
   48241: out<=1;
   48242: out<=1;
   48243: out<=1;
   48244: out<=0;
   48245: out<=1;
   48246: out<=1;
   48247: out<=0;
   48248: out<=1;
   48249: out<=0;
   48250: out<=1;
   48251: out<=0;
   48252: out<=0;
   48253: out<=0;
   48254: out<=1;
   48255: out<=1;
   48256: out<=0;
   48257: out<=0;
   48258: out<=0;
   48259: out<=0;
   48260: out<=1;
   48261: out<=0;
   48262: out<=0;
   48263: out<=1;
   48264: out<=0;
   48265: out<=1;
   48266: out<=0;
   48267: out<=1;
   48268: out<=1;
   48269: out<=1;
   48270: out<=0;
   48271: out<=0;
   48272: out<=1;
   48273: out<=1;
   48274: out<=1;
   48275: out<=1;
   48276: out<=0;
   48277: out<=1;
   48278: out<=1;
   48279: out<=0;
   48280: out<=1;
   48281: out<=0;
   48282: out<=1;
   48283: out<=0;
   48284: out<=0;
   48285: out<=0;
   48286: out<=1;
   48287: out<=1;
   48288: out<=1;
   48289: out<=1;
   48290: out<=1;
   48291: out<=1;
   48292: out<=0;
   48293: out<=1;
   48294: out<=1;
   48295: out<=0;
   48296: out<=1;
   48297: out<=0;
   48298: out<=1;
   48299: out<=0;
   48300: out<=0;
   48301: out<=0;
   48302: out<=1;
   48303: out<=1;
   48304: out<=0;
   48305: out<=0;
   48306: out<=0;
   48307: out<=0;
   48308: out<=1;
   48309: out<=0;
   48310: out<=0;
   48311: out<=1;
   48312: out<=0;
   48313: out<=1;
   48314: out<=0;
   48315: out<=1;
   48316: out<=1;
   48317: out<=1;
   48318: out<=0;
   48319: out<=0;
   48320: out<=1;
   48321: out<=1;
   48322: out<=1;
   48323: out<=1;
   48324: out<=0;
   48325: out<=1;
   48326: out<=1;
   48327: out<=0;
   48328: out<=1;
   48329: out<=0;
   48330: out<=1;
   48331: out<=0;
   48332: out<=0;
   48333: out<=0;
   48334: out<=1;
   48335: out<=1;
   48336: out<=1;
   48337: out<=1;
   48338: out<=1;
   48339: out<=1;
   48340: out<=0;
   48341: out<=1;
   48342: out<=1;
   48343: out<=0;
   48344: out<=1;
   48345: out<=0;
   48346: out<=1;
   48347: out<=0;
   48348: out<=0;
   48349: out<=0;
   48350: out<=1;
   48351: out<=1;
   48352: out<=1;
   48353: out<=1;
   48354: out<=1;
   48355: out<=1;
   48356: out<=0;
   48357: out<=1;
   48358: out<=1;
   48359: out<=0;
   48360: out<=1;
   48361: out<=0;
   48362: out<=1;
   48363: out<=0;
   48364: out<=0;
   48365: out<=0;
   48366: out<=1;
   48367: out<=1;
   48368: out<=1;
   48369: out<=1;
   48370: out<=1;
   48371: out<=1;
   48372: out<=0;
   48373: out<=1;
   48374: out<=1;
   48375: out<=0;
   48376: out<=1;
   48377: out<=0;
   48378: out<=1;
   48379: out<=0;
   48380: out<=0;
   48381: out<=0;
   48382: out<=1;
   48383: out<=1;
   48384: out<=1;
   48385: out<=0;
   48386: out<=0;
   48387: out<=1;
   48388: out<=1;
   48389: out<=1;
   48390: out<=1;
   48391: out<=1;
   48392: out<=0;
   48393: out<=0;
   48394: out<=1;
   48395: out<=1;
   48396: out<=0;
   48397: out<=1;
   48398: out<=0;
   48399: out<=1;
   48400: out<=0;
   48401: out<=1;
   48402: out<=1;
   48403: out<=0;
   48404: out<=0;
   48405: out<=0;
   48406: out<=0;
   48407: out<=0;
   48408: out<=1;
   48409: out<=1;
   48410: out<=0;
   48411: out<=0;
   48412: out<=1;
   48413: out<=0;
   48414: out<=1;
   48415: out<=0;
   48416: out<=1;
   48417: out<=0;
   48418: out<=0;
   48419: out<=1;
   48420: out<=1;
   48421: out<=1;
   48422: out<=1;
   48423: out<=1;
   48424: out<=0;
   48425: out<=0;
   48426: out<=1;
   48427: out<=1;
   48428: out<=0;
   48429: out<=1;
   48430: out<=0;
   48431: out<=1;
   48432: out<=0;
   48433: out<=1;
   48434: out<=1;
   48435: out<=0;
   48436: out<=0;
   48437: out<=0;
   48438: out<=0;
   48439: out<=0;
   48440: out<=1;
   48441: out<=1;
   48442: out<=0;
   48443: out<=0;
   48444: out<=1;
   48445: out<=0;
   48446: out<=1;
   48447: out<=0;
   48448: out<=0;
   48449: out<=1;
   48450: out<=1;
   48451: out<=0;
   48452: out<=0;
   48453: out<=0;
   48454: out<=0;
   48455: out<=0;
   48456: out<=1;
   48457: out<=1;
   48458: out<=0;
   48459: out<=0;
   48460: out<=1;
   48461: out<=0;
   48462: out<=1;
   48463: out<=0;
   48464: out<=0;
   48465: out<=1;
   48466: out<=1;
   48467: out<=0;
   48468: out<=0;
   48469: out<=0;
   48470: out<=0;
   48471: out<=0;
   48472: out<=1;
   48473: out<=1;
   48474: out<=0;
   48475: out<=0;
   48476: out<=1;
   48477: out<=0;
   48478: out<=1;
   48479: out<=0;
   48480: out<=1;
   48481: out<=0;
   48482: out<=0;
   48483: out<=1;
   48484: out<=1;
   48485: out<=1;
   48486: out<=1;
   48487: out<=1;
   48488: out<=0;
   48489: out<=0;
   48490: out<=1;
   48491: out<=1;
   48492: out<=0;
   48493: out<=1;
   48494: out<=0;
   48495: out<=1;
   48496: out<=1;
   48497: out<=0;
   48498: out<=0;
   48499: out<=1;
   48500: out<=1;
   48501: out<=1;
   48502: out<=1;
   48503: out<=1;
   48504: out<=0;
   48505: out<=0;
   48506: out<=1;
   48507: out<=1;
   48508: out<=0;
   48509: out<=1;
   48510: out<=0;
   48511: out<=1;
   48512: out<=0;
   48513: out<=1;
   48514: out<=1;
   48515: out<=0;
   48516: out<=0;
   48517: out<=0;
   48518: out<=0;
   48519: out<=0;
   48520: out<=1;
   48521: out<=1;
   48522: out<=0;
   48523: out<=0;
   48524: out<=1;
   48525: out<=0;
   48526: out<=1;
   48527: out<=0;
   48528: out<=0;
   48529: out<=1;
   48530: out<=1;
   48531: out<=0;
   48532: out<=0;
   48533: out<=0;
   48534: out<=0;
   48535: out<=0;
   48536: out<=1;
   48537: out<=1;
   48538: out<=0;
   48539: out<=0;
   48540: out<=1;
   48541: out<=0;
   48542: out<=1;
   48543: out<=0;
   48544: out<=0;
   48545: out<=1;
   48546: out<=1;
   48547: out<=0;
   48548: out<=0;
   48549: out<=0;
   48550: out<=0;
   48551: out<=0;
   48552: out<=1;
   48553: out<=1;
   48554: out<=0;
   48555: out<=0;
   48556: out<=1;
   48557: out<=0;
   48558: out<=1;
   48559: out<=0;
   48560: out<=0;
   48561: out<=1;
   48562: out<=1;
   48563: out<=0;
   48564: out<=0;
   48565: out<=0;
   48566: out<=0;
   48567: out<=0;
   48568: out<=1;
   48569: out<=1;
   48570: out<=0;
   48571: out<=0;
   48572: out<=1;
   48573: out<=0;
   48574: out<=1;
   48575: out<=0;
   48576: out<=1;
   48577: out<=0;
   48578: out<=0;
   48579: out<=1;
   48580: out<=1;
   48581: out<=1;
   48582: out<=1;
   48583: out<=1;
   48584: out<=0;
   48585: out<=0;
   48586: out<=1;
   48587: out<=1;
   48588: out<=0;
   48589: out<=1;
   48590: out<=0;
   48591: out<=1;
   48592: out<=0;
   48593: out<=1;
   48594: out<=1;
   48595: out<=0;
   48596: out<=0;
   48597: out<=0;
   48598: out<=0;
   48599: out<=0;
   48600: out<=1;
   48601: out<=1;
   48602: out<=0;
   48603: out<=0;
   48604: out<=1;
   48605: out<=0;
   48606: out<=1;
   48607: out<=0;
   48608: out<=0;
   48609: out<=1;
   48610: out<=1;
   48611: out<=0;
   48612: out<=0;
   48613: out<=0;
   48614: out<=0;
   48615: out<=0;
   48616: out<=1;
   48617: out<=1;
   48618: out<=0;
   48619: out<=0;
   48620: out<=1;
   48621: out<=0;
   48622: out<=1;
   48623: out<=0;
   48624: out<=1;
   48625: out<=0;
   48626: out<=0;
   48627: out<=1;
   48628: out<=1;
   48629: out<=1;
   48630: out<=1;
   48631: out<=1;
   48632: out<=0;
   48633: out<=0;
   48634: out<=1;
   48635: out<=1;
   48636: out<=0;
   48637: out<=1;
   48638: out<=0;
   48639: out<=1;
   48640: out<=0;
   48641: out<=1;
   48642: out<=0;
   48643: out<=1;
   48644: out<=0;
   48645: out<=0;
   48646: out<=1;
   48647: out<=1;
   48648: out<=0;
   48649: out<=0;
   48650: out<=0;
   48651: out<=0;
   48652: out<=0;
   48653: out<=1;
   48654: out<=1;
   48655: out<=0;
   48656: out<=1;
   48657: out<=0;
   48658: out<=1;
   48659: out<=0;
   48660: out<=1;
   48661: out<=1;
   48662: out<=0;
   48663: out<=0;
   48664: out<=1;
   48665: out<=1;
   48666: out<=1;
   48667: out<=1;
   48668: out<=1;
   48669: out<=0;
   48670: out<=0;
   48671: out<=1;
   48672: out<=1;
   48673: out<=0;
   48674: out<=1;
   48675: out<=0;
   48676: out<=1;
   48677: out<=1;
   48678: out<=0;
   48679: out<=0;
   48680: out<=1;
   48681: out<=1;
   48682: out<=1;
   48683: out<=1;
   48684: out<=1;
   48685: out<=0;
   48686: out<=0;
   48687: out<=1;
   48688: out<=0;
   48689: out<=1;
   48690: out<=0;
   48691: out<=1;
   48692: out<=0;
   48693: out<=0;
   48694: out<=1;
   48695: out<=1;
   48696: out<=0;
   48697: out<=0;
   48698: out<=0;
   48699: out<=0;
   48700: out<=0;
   48701: out<=1;
   48702: out<=1;
   48703: out<=0;
   48704: out<=1;
   48705: out<=0;
   48706: out<=1;
   48707: out<=0;
   48708: out<=1;
   48709: out<=1;
   48710: out<=0;
   48711: out<=0;
   48712: out<=1;
   48713: out<=1;
   48714: out<=1;
   48715: out<=1;
   48716: out<=1;
   48717: out<=0;
   48718: out<=0;
   48719: out<=1;
   48720: out<=1;
   48721: out<=0;
   48722: out<=1;
   48723: out<=0;
   48724: out<=1;
   48725: out<=1;
   48726: out<=0;
   48727: out<=0;
   48728: out<=1;
   48729: out<=1;
   48730: out<=1;
   48731: out<=1;
   48732: out<=1;
   48733: out<=0;
   48734: out<=0;
   48735: out<=1;
   48736: out<=1;
   48737: out<=0;
   48738: out<=1;
   48739: out<=0;
   48740: out<=1;
   48741: out<=1;
   48742: out<=0;
   48743: out<=0;
   48744: out<=1;
   48745: out<=1;
   48746: out<=1;
   48747: out<=1;
   48748: out<=1;
   48749: out<=0;
   48750: out<=0;
   48751: out<=1;
   48752: out<=1;
   48753: out<=0;
   48754: out<=1;
   48755: out<=0;
   48756: out<=1;
   48757: out<=1;
   48758: out<=0;
   48759: out<=0;
   48760: out<=1;
   48761: out<=1;
   48762: out<=1;
   48763: out<=1;
   48764: out<=1;
   48765: out<=0;
   48766: out<=0;
   48767: out<=1;
   48768: out<=1;
   48769: out<=0;
   48770: out<=1;
   48771: out<=0;
   48772: out<=1;
   48773: out<=1;
   48774: out<=0;
   48775: out<=0;
   48776: out<=1;
   48777: out<=1;
   48778: out<=1;
   48779: out<=1;
   48780: out<=1;
   48781: out<=0;
   48782: out<=0;
   48783: out<=1;
   48784: out<=1;
   48785: out<=0;
   48786: out<=1;
   48787: out<=0;
   48788: out<=1;
   48789: out<=1;
   48790: out<=0;
   48791: out<=0;
   48792: out<=1;
   48793: out<=1;
   48794: out<=1;
   48795: out<=1;
   48796: out<=1;
   48797: out<=0;
   48798: out<=0;
   48799: out<=1;
   48800: out<=0;
   48801: out<=1;
   48802: out<=0;
   48803: out<=1;
   48804: out<=0;
   48805: out<=0;
   48806: out<=1;
   48807: out<=1;
   48808: out<=0;
   48809: out<=0;
   48810: out<=0;
   48811: out<=0;
   48812: out<=0;
   48813: out<=1;
   48814: out<=1;
   48815: out<=0;
   48816: out<=0;
   48817: out<=1;
   48818: out<=0;
   48819: out<=1;
   48820: out<=0;
   48821: out<=0;
   48822: out<=1;
   48823: out<=1;
   48824: out<=0;
   48825: out<=0;
   48826: out<=0;
   48827: out<=0;
   48828: out<=0;
   48829: out<=1;
   48830: out<=1;
   48831: out<=0;
   48832: out<=0;
   48833: out<=1;
   48834: out<=0;
   48835: out<=1;
   48836: out<=0;
   48837: out<=0;
   48838: out<=1;
   48839: out<=1;
   48840: out<=0;
   48841: out<=0;
   48842: out<=0;
   48843: out<=0;
   48844: out<=0;
   48845: out<=1;
   48846: out<=1;
   48847: out<=0;
   48848: out<=1;
   48849: out<=0;
   48850: out<=1;
   48851: out<=0;
   48852: out<=1;
   48853: out<=1;
   48854: out<=0;
   48855: out<=0;
   48856: out<=1;
   48857: out<=1;
   48858: out<=1;
   48859: out<=1;
   48860: out<=1;
   48861: out<=0;
   48862: out<=0;
   48863: out<=1;
   48864: out<=0;
   48865: out<=1;
   48866: out<=0;
   48867: out<=1;
   48868: out<=0;
   48869: out<=0;
   48870: out<=1;
   48871: out<=1;
   48872: out<=0;
   48873: out<=0;
   48874: out<=0;
   48875: out<=0;
   48876: out<=0;
   48877: out<=1;
   48878: out<=1;
   48879: out<=0;
   48880: out<=1;
   48881: out<=0;
   48882: out<=1;
   48883: out<=0;
   48884: out<=1;
   48885: out<=1;
   48886: out<=0;
   48887: out<=0;
   48888: out<=1;
   48889: out<=1;
   48890: out<=1;
   48891: out<=1;
   48892: out<=1;
   48893: out<=0;
   48894: out<=0;
   48895: out<=1;
   48896: out<=0;
   48897: out<=0;
   48898: out<=1;
   48899: out<=1;
   48900: out<=1;
   48901: out<=0;
   48902: out<=1;
   48903: out<=0;
   48904: out<=1;
   48905: out<=0;
   48906: out<=0;
   48907: out<=1;
   48908: out<=0;
   48909: out<=0;
   48910: out<=0;
   48911: out<=0;
   48912: out<=0;
   48913: out<=0;
   48914: out<=1;
   48915: out<=1;
   48916: out<=1;
   48917: out<=0;
   48918: out<=1;
   48919: out<=0;
   48920: out<=1;
   48921: out<=0;
   48922: out<=0;
   48923: out<=1;
   48924: out<=0;
   48925: out<=0;
   48926: out<=0;
   48927: out<=0;
   48928: out<=0;
   48929: out<=0;
   48930: out<=1;
   48931: out<=1;
   48932: out<=1;
   48933: out<=0;
   48934: out<=1;
   48935: out<=0;
   48936: out<=1;
   48937: out<=0;
   48938: out<=0;
   48939: out<=1;
   48940: out<=0;
   48941: out<=0;
   48942: out<=0;
   48943: out<=0;
   48944: out<=0;
   48945: out<=0;
   48946: out<=1;
   48947: out<=1;
   48948: out<=1;
   48949: out<=0;
   48950: out<=1;
   48951: out<=0;
   48952: out<=1;
   48953: out<=0;
   48954: out<=0;
   48955: out<=1;
   48956: out<=0;
   48957: out<=0;
   48958: out<=0;
   48959: out<=0;
   48960: out<=1;
   48961: out<=1;
   48962: out<=0;
   48963: out<=0;
   48964: out<=0;
   48965: out<=1;
   48966: out<=0;
   48967: out<=1;
   48968: out<=0;
   48969: out<=1;
   48970: out<=1;
   48971: out<=0;
   48972: out<=1;
   48973: out<=1;
   48974: out<=1;
   48975: out<=1;
   48976: out<=0;
   48977: out<=0;
   48978: out<=1;
   48979: out<=1;
   48980: out<=1;
   48981: out<=0;
   48982: out<=1;
   48983: out<=0;
   48984: out<=1;
   48985: out<=0;
   48986: out<=0;
   48987: out<=1;
   48988: out<=0;
   48989: out<=0;
   48990: out<=0;
   48991: out<=0;
   48992: out<=0;
   48993: out<=0;
   48994: out<=1;
   48995: out<=1;
   48996: out<=1;
   48997: out<=0;
   48998: out<=1;
   48999: out<=0;
   49000: out<=1;
   49001: out<=0;
   49002: out<=0;
   49003: out<=1;
   49004: out<=0;
   49005: out<=0;
   49006: out<=0;
   49007: out<=0;
   49008: out<=1;
   49009: out<=1;
   49010: out<=0;
   49011: out<=0;
   49012: out<=0;
   49013: out<=1;
   49014: out<=0;
   49015: out<=1;
   49016: out<=0;
   49017: out<=1;
   49018: out<=1;
   49019: out<=0;
   49020: out<=1;
   49021: out<=1;
   49022: out<=1;
   49023: out<=1;
   49024: out<=1;
   49025: out<=1;
   49026: out<=0;
   49027: out<=0;
   49028: out<=0;
   49029: out<=1;
   49030: out<=0;
   49031: out<=1;
   49032: out<=0;
   49033: out<=1;
   49034: out<=1;
   49035: out<=0;
   49036: out<=1;
   49037: out<=1;
   49038: out<=1;
   49039: out<=1;
   49040: out<=0;
   49041: out<=0;
   49042: out<=1;
   49043: out<=1;
   49044: out<=1;
   49045: out<=0;
   49046: out<=1;
   49047: out<=0;
   49048: out<=1;
   49049: out<=0;
   49050: out<=0;
   49051: out<=1;
   49052: out<=0;
   49053: out<=0;
   49054: out<=0;
   49055: out<=0;
   49056: out<=1;
   49057: out<=1;
   49058: out<=0;
   49059: out<=0;
   49060: out<=0;
   49061: out<=1;
   49062: out<=0;
   49063: out<=1;
   49064: out<=0;
   49065: out<=1;
   49066: out<=1;
   49067: out<=0;
   49068: out<=1;
   49069: out<=1;
   49070: out<=1;
   49071: out<=1;
   49072: out<=0;
   49073: out<=0;
   49074: out<=1;
   49075: out<=1;
   49076: out<=1;
   49077: out<=0;
   49078: out<=1;
   49079: out<=0;
   49080: out<=1;
   49081: out<=0;
   49082: out<=0;
   49083: out<=1;
   49084: out<=0;
   49085: out<=0;
   49086: out<=0;
   49087: out<=0;
   49088: out<=0;
   49089: out<=0;
   49090: out<=1;
   49091: out<=1;
   49092: out<=1;
   49093: out<=0;
   49094: out<=1;
   49095: out<=0;
   49096: out<=1;
   49097: out<=0;
   49098: out<=0;
   49099: out<=1;
   49100: out<=0;
   49101: out<=0;
   49102: out<=0;
   49103: out<=0;
   49104: out<=0;
   49105: out<=0;
   49106: out<=1;
   49107: out<=1;
   49108: out<=1;
   49109: out<=0;
   49110: out<=1;
   49111: out<=0;
   49112: out<=1;
   49113: out<=0;
   49114: out<=0;
   49115: out<=1;
   49116: out<=0;
   49117: out<=0;
   49118: out<=0;
   49119: out<=0;
   49120: out<=1;
   49121: out<=1;
   49122: out<=0;
   49123: out<=0;
   49124: out<=0;
   49125: out<=1;
   49126: out<=0;
   49127: out<=1;
   49128: out<=0;
   49129: out<=1;
   49130: out<=1;
   49131: out<=0;
   49132: out<=1;
   49133: out<=1;
   49134: out<=1;
   49135: out<=1;
   49136: out<=1;
   49137: out<=1;
   49138: out<=0;
   49139: out<=0;
   49140: out<=0;
   49141: out<=1;
   49142: out<=0;
   49143: out<=1;
   49144: out<=0;
   49145: out<=1;
   49146: out<=1;
   49147: out<=0;
   49148: out<=1;
   49149: out<=1;
   49150: out<=1;
   49151: out<=1;
   49152: out<=0;
   49153: out<=0;
   49154: out<=0;
   49155: out<=0;
   49156: out<=1;
   49157: out<=0;
   49158: out<=0;
   49159: out<=1;
   49160: out<=0;
   49161: out<=1;
   49162: out<=0;
   49163: out<=1;
   49164: out<=1;
   49165: out<=1;
   49166: out<=0;
   49167: out<=0;
   49168: out<=1;
   49169: out<=1;
   49170: out<=1;
   49171: out<=1;
   49172: out<=0;
   49173: out<=1;
   49174: out<=1;
   49175: out<=0;
   49176: out<=1;
   49177: out<=0;
   49178: out<=1;
   49179: out<=0;
   49180: out<=0;
   49181: out<=0;
   49182: out<=1;
   49183: out<=1;
   49184: out<=1;
   49185: out<=1;
   49186: out<=1;
   49187: out<=1;
   49188: out<=0;
   49189: out<=1;
   49190: out<=1;
   49191: out<=0;
   49192: out<=1;
   49193: out<=0;
   49194: out<=1;
   49195: out<=0;
   49196: out<=0;
   49197: out<=0;
   49198: out<=1;
   49199: out<=1;
   49200: out<=0;
   49201: out<=0;
   49202: out<=0;
   49203: out<=0;
   49204: out<=1;
   49205: out<=0;
   49206: out<=0;
   49207: out<=1;
   49208: out<=0;
   49209: out<=1;
   49210: out<=0;
   49211: out<=1;
   49212: out<=1;
   49213: out<=1;
   49214: out<=0;
   49215: out<=0;
   49216: out<=1;
   49217: out<=1;
   49218: out<=1;
   49219: out<=1;
   49220: out<=0;
   49221: out<=1;
   49222: out<=1;
   49223: out<=0;
   49224: out<=1;
   49225: out<=0;
   49226: out<=1;
   49227: out<=0;
   49228: out<=0;
   49229: out<=0;
   49230: out<=1;
   49231: out<=1;
   49232: out<=1;
   49233: out<=1;
   49234: out<=1;
   49235: out<=1;
   49236: out<=0;
   49237: out<=1;
   49238: out<=1;
   49239: out<=0;
   49240: out<=1;
   49241: out<=0;
   49242: out<=1;
   49243: out<=0;
   49244: out<=0;
   49245: out<=0;
   49246: out<=1;
   49247: out<=1;
   49248: out<=1;
   49249: out<=1;
   49250: out<=1;
   49251: out<=1;
   49252: out<=0;
   49253: out<=1;
   49254: out<=1;
   49255: out<=0;
   49256: out<=1;
   49257: out<=0;
   49258: out<=1;
   49259: out<=0;
   49260: out<=0;
   49261: out<=0;
   49262: out<=1;
   49263: out<=1;
   49264: out<=1;
   49265: out<=1;
   49266: out<=1;
   49267: out<=1;
   49268: out<=0;
   49269: out<=1;
   49270: out<=1;
   49271: out<=0;
   49272: out<=1;
   49273: out<=0;
   49274: out<=1;
   49275: out<=0;
   49276: out<=0;
   49277: out<=0;
   49278: out<=1;
   49279: out<=1;
   49280: out<=0;
   49281: out<=0;
   49282: out<=0;
   49283: out<=0;
   49284: out<=1;
   49285: out<=0;
   49286: out<=0;
   49287: out<=1;
   49288: out<=0;
   49289: out<=1;
   49290: out<=0;
   49291: out<=1;
   49292: out<=1;
   49293: out<=1;
   49294: out<=0;
   49295: out<=0;
   49296: out<=0;
   49297: out<=0;
   49298: out<=0;
   49299: out<=0;
   49300: out<=1;
   49301: out<=0;
   49302: out<=0;
   49303: out<=1;
   49304: out<=0;
   49305: out<=1;
   49306: out<=0;
   49307: out<=1;
   49308: out<=1;
   49309: out<=1;
   49310: out<=0;
   49311: out<=0;
   49312: out<=1;
   49313: out<=1;
   49314: out<=1;
   49315: out<=1;
   49316: out<=0;
   49317: out<=1;
   49318: out<=1;
   49319: out<=0;
   49320: out<=1;
   49321: out<=0;
   49322: out<=1;
   49323: out<=0;
   49324: out<=0;
   49325: out<=0;
   49326: out<=1;
   49327: out<=1;
   49328: out<=1;
   49329: out<=1;
   49330: out<=1;
   49331: out<=1;
   49332: out<=0;
   49333: out<=1;
   49334: out<=1;
   49335: out<=0;
   49336: out<=1;
   49337: out<=0;
   49338: out<=1;
   49339: out<=0;
   49340: out<=0;
   49341: out<=0;
   49342: out<=1;
   49343: out<=1;
   49344: out<=1;
   49345: out<=1;
   49346: out<=1;
   49347: out<=1;
   49348: out<=0;
   49349: out<=1;
   49350: out<=1;
   49351: out<=0;
   49352: out<=1;
   49353: out<=0;
   49354: out<=1;
   49355: out<=0;
   49356: out<=0;
   49357: out<=0;
   49358: out<=1;
   49359: out<=1;
   49360: out<=0;
   49361: out<=0;
   49362: out<=0;
   49363: out<=0;
   49364: out<=1;
   49365: out<=0;
   49366: out<=0;
   49367: out<=1;
   49368: out<=0;
   49369: out<=1;
   49370: out<=0;
   49371: out<=1;
   49372: out<=1;
   49373: out<=1;
   49374: out<=0;
   49375: out<=0;
   49376: out<=1;
   49377: out<=1;
   49378: out<=1;
   49379: out<=1;
   49380: out<=0;
   49381: out<=1;
   49382: out<=1;
   49383: out<=0;
   49384: out<=1;
   49385: out<=0;
   49386: out<=1;
   49387: out<=0;
   49388: out<=0;
   49389: out<=0;
   49390: out<=1;
   49391: out<=1;
   49392: out<=0;
   49393: out<=0;
   49394: out<=0;
   49395: out<=0;
   49396: out<=1;
   49397: out<=0;
   49398: out<=0;
   49399: out<=1;
   49400: out<=0;
   49401: out<=1;
   49402: out<=0;
   49403: out<=1;
   49404: out<=1;
   49405: out<=1;
   49406: out<=0;
   49407: out<=0;
   49408: out<=0;
   49409: out<=1;
   49410: out<=1;
   49411: out<=0;
   49412: out<=0;
   49413: out<=0;
   49414: out<=0;
   49415: out<=0;
   49416: out<=1;
   49417: out<=1;
   49418: out<=0;
   49419: out<=0;
   49420: out<=1;
   49421: out<=0;
   49422: out<=1;
   49423: out<=0;
   49424: out<=0;
   49425: out<=1;
   49426: out<=1;
   49427: out<=0;
   49428: out<=0;
   49429: out<=0;
   49430: out<=0;
   49431: out<=0;
   49432: out<=1;
   49433: out<=1;
   49434: out<=0;
   49435: out<=0;
   49436: out<=1;
   49437: out<=0;
   49438: out<=1;
   49439: out<=0;
   49440: out<=0;
   49441: out<=1;
   49442: out<=1;
   49443: out<=0;
   49444: out<=0;
   49445: out<=0;
   49446: out<=0;
   49447: out<=0;
   49448: out<=1;
   49449: out<=1;
   49450: out<=0;
   49451: out<=0;
   49452: out<=1;
   49453: out<=0;
   49454: out<=1;
   49455: out<=0;
   49456: out<=0;
   49457: out<=1;
   49458: out<=1;
   49459: out<=0;
   49460: out<=0;
   49461: out<=0;
   49462: out<=0;
   49463: out<=0;
   49464: out<=1;
   49465: out<=1;
   49466: out<=0;
   49467: out<=0;
   49468: out<=1;
   49469: out<=0;
   49470: out<=1;
   49471: out<=0;
   49472: out<=1;
   49473: out<=0;
   49474: out<=0;
   49475: out<=1;
   49476: out<=1;
   49477: out<=1;
   49478: out<=1;
   49479: out<=1;
   49480: out<=0;
   49481: out<=0;
   49482: out<=1;
   49483: out<=1;
   49484: out<=0;
   49485: out<=1;
   49486: out<=0;
   49487: out<=1;
   49488: out<=0;
   49489: out<=1;
   49490: out<=1;
   49491: out<=0;
   49492: out<=0;
   49493: out<=0;
   49494: out<=0;
   49495: out<=0;
   49496: out<=1;
   49497: out<=1;
   49498: out<=0;
   49499: out<=0;
   49500: out<=1;
   49501: out<=0;
   49502: out<=1;
   49503: out<=0;
   49504: out<=0;
   49505: out<=1;
   49506: out<=1;
   49507: out<=0;
   49508: out<=0;
   49509: out<=0;
   49510: out<=0;
   49511: out<=0;
   49512: out<=1;
   49513: out<=1;
   49514: out<=0;
   49515: out<=0;
   49516: out<=1;
   49517: out<=0;
   49518: out<=1;
   49519: out<=0;
   49520: out<=1;
   49521: out<=0;
   49522: out<=0;
   49523: out<=1;
   49524: out<=1;
   49525: out<=1;
   49526: out<=1;
   49527: out<=1;
   49528: out<=0;
   49529: out<=0;
   49530: out<=1;
   49531: out<=1;
   49532: out<=0;
   49533: out<=1;
   49534: out<=0;
   49535: out<=1;
   49536: out<=0;
   49537: out<=1;
   49538: out<=1;
   49539: out<=0;
   49540: out<=0;
   49541: out<=0;
   49542: out<=0;
   49543: out<=0;
   49544: out<=1;
   49545: out<=1;
   49546: out<=0;
   49547: out<=0;
   49548: out<=1;
   49549: out<=0;
   49550: out<=1;
   49551: out<=0;
   49552: out<=1;
   49553: out<=0;
   49554: out<=0;
   49555: out<=1;
   49556: out<=1;
   49557: out<=1;
   49558: out<=1;
   49559: out<=1;
   49560: out<=0;
   49561: out<=0;
   49562: out<=1;
   49563: out<=1;
   49564: out<=0;
   49565: out<=1;
   49566: out<=0;
   49567: out<=1;
   49568: out<=0;
   49569: out<=1;
   49570: out<=1;
   49571: out<=0;
   49572: out<=0;
   49573: out<=0;
   49574: out<=0;
   49575: out<=0;
   49576: out<=1;
   49577: out<=1;
   49578: out<=0;
   49579: out<=0;
   49580: out<=1;
   49581: out<=0;
   49582: out<=1;
   49583: out<=0;
   49584: out<=1;
   49585: out<=0;
   49586: out<=0;
   49587: out<=1;
   49588: out<=1;
   49589: out<=1;
   49590: out<=1;
   49591: out<=1;
   49592: out<=0;
   49593: out<=0;
   49594: out<=1;
   49595: out<=1;
   49596: out<=0;
   49597: out<=1;
   49598: out<=0;
   49599: out<=1;
   49600: out<=1;
   49601: out<=0;
   49602: out<=0;
   49603: out<=1;
   49604: out<=1;
   49605: out<=1;
   49606: out<=1;
   49607: out<=1;
   49608: out<=0;
   49609: out<=0;
   49610: out<=1;
   49611: out<=1;
   49612: out<=0;
   49613: out<=1;
   49614: out<=0;
   49615: out<=1;
   49616: out<=1;
   49617: out<=0;
   49618: out<=0;
   49619: out<=1;
   49620: out<=1;
   49621: out<=1;
   49622: out<=1;
   49623: out<=1;
   49624: out<=0;
   49625: out<=0;
   49626: out<=1;
   49627: out<=1;
   49628: out<=0;
   49629: out<=1;
   49630: out<=0;
   49631: out<=1;
   49632: out<=0;
   49633: out<=1;
   49634: out<=1;
   49635: out<=0;
   49636: out<=0;
   49637: out<=0;
   49638: out<=0;
   49639: out<=0;
   49640: out<=1;
   49641: out<=1;
   49642: out<=0;
   49643: out<=0;
   49644: out<=1;
   49645: out<=0;
   49646: out<=1;
   49647: out<=0;
   49648: out<=0;
   49649: out<=1;
   49650: out<=1;
   49651: out<=0;
   49652: out<=0;
   49653: out<=0;
   49654: out<=0;
   49655: out<=0;
   49656: out<=1;
   49657: out<=1;
   49658: out<=0;
   49659: out<=0;
   49660: out<=1;
   49661: out<=0;
   49662: out<=1;
   49663: out<=0;
   49664: out<=0;
   49665: out<=1;
   49666: out<=0;
   49667: out<=1;
   49668: out<=0;
   49669: out<=0;
   49670: out<=1;
   49671: out<=1;
   49672: out<=0;
   49673: out<=0;
   49674: out<=0;
   49675: out<=0;
   49676: out<=0;
   49677: out<=1;
   49678: out<=1;
   49679: out<=0;
   49680: out<=0;
   49681: out<=1;
   49682: out<=0;
   49683: out<=1;
   49684: out<=0;
   49685: out<=0;
   49686: out<=1;
   49687: out<=1;
   49688: out<=0;
   49689: out<=0;
   49690: out<=0;
   49691: out<=0;
   49692: out<=0;
   49693: out<=1;
   49694: out<=1;
   49695: out<=0;
   49696: out<=1;
   49697: out<=0;
   49698: out<=1;
   49699: out<=0;
   49700: out<=1;
   49701: out<=1;
   49702: out<=0;
   49703: out<=0;
   49704: out<=1;
   49705: out<=1;
   49706: out<=1;
   49707: out<=1;
   49708: out<=1;
   49709: out<=0;
   49710: out<=0;
   49711: out<=1;
   49712: out<=1;
   49713: out<=0;
   49714: out<=1;
   49715: out<=0;
   49716: out<=1;
   49717: out<=1;
   49718: out<=0;
   49719: out<=0;
   49720: out<=1;
   49721: out<=1;
   49722: out<=1;
   49723: out<=1;
   49724: out<=1;
   49725: out<=0;
   49726: out<=0;
   49727: out<=1;
   49728: out<=1;
   49729: out<=0;
   49730: out<=1;
   49731: out<=0;
   49732: out<=1;
   49733: out<=1;
   49734: out<=0;
   49735: out<=0;
   49736: out<=1;
   49737: out<=1;
   49738: out<=1;
   49739: out<=1;
   49740: out<=1;
   49741: out<=0;
   49742: out<=0;
   49743: out<=1;
   49744: out<=0;
   49745: out<=1;
   49746: out<=0;
   49747: out<=1;
   49748: out<=0;
   49749: out<=0;
   49750: out<=1;
   49751: out<=1;
   49752: out<=0;
   49753: out<=0;
   49754: out<=0;
   49755: out<=0;
   49756: out<=0;
   49757: out<=1;
   49758: out<=1;
   49759: out<=0;
   49760: out<=1;
   49761: out<=0;
   49762: out<=1;
   49763: out<=0;
   49764: out<=1;
   49765: out<=1;
   49766: out<=0;
   49767: out<=0;
   49768: out<=1;
   49769: out<=1;
   49770: out<=1;
   49771: out<=1;
   49772: out<=1;
   49773: out<=0;
   49774: out<=0;
   49775: out<=1;
   49776: out<=0;
   49777: out<=1;
   49778: out<=0;
   49779: out<=1;
   49780: out<=0;
   49781: out<=0;
   49782: out<=1;
   49783: out<=1;
   49784: out<=0;
   49785: out<=0;
   49786: out<=0;
   49787: out<=0;
   49788: out<=0;
   49789: out<=1;
   49790: out<=1;
   49791: out<=0;
   49792: out<=0;
   49793: out<=1;
   49794: out<=0;
   49795: out<=1;
   49796: out<=0;
   49797: out<=0;
   49798: out<=1;
   49799: out<=1;
   49800: out<=0;
   49801: out<=0;
   49802: out<=0;
   49803: out<=0;
   49804: out<=0;
   49805: out<=1;
   49806: out<=1;
   49807: out<=0;
   49808: out<=1;
   49809: out<=0;
   49810: out<=1;
   49811: out<=0;
   49812: out<=1;
   49813: out<=1;
   49814: out<=0;
   49815: out<=0;
   49816: out<=1;
   49817: out<=1;
   49818: out<=1;
   49819: out<=1;
   49820: out<=1;
   49821: out<=0;
   49822: out<=0;
   49823: out<=1;
   49824: out<=1;
   49825: out<=0;
   49826: out<=1;
   49827: out<=0;
   49828: out<=1;
   49829: out<=1;
   49830: out<=0;
   49831: out<=0;
   49832: out<=1;
   49833: out<=1;
   49834: out<=1;
   49835: out<=1;
   49836: out<=1;
   49837: out<=0;
   49838: out<=0;
   49839: out<=1;
   49840: out<=0;
   49841: out<=1;
   49842: out<=0;
   49843: out<=1;
   49844: out<=0;
   49845: out<=0;
   49846: out<=1;
   49847: out<=1;
   49848: out<=0;
   49849: out<=0;
   49850: out<=0;
   49851: out<=0;
   49852: out<=0;
   49853: out<=1;
   49854: out<=1;
   49855: out<=0;
   49856: out<=1;
   49857: out<=0;
   49858: out<=1;
   49859: out<=0;
   49860: out<=1;
   49861: out<=1;
   49862: out<=0;
   49863: out<=0;
   49864: out<=1;
   49865: out<=1;
   49866: out<=1;
   49867: out<=1;
   49868: out<=1;
   49869: out<=0;
   49870: out<=0;
   49871: out<=1;
   49872: out<=1;
   49873: out<=0;
   49874: out<=1;
   49875: out<=0;
   49876: out<=1;
   49877: out<=1;
   49878: out<=0;
   49879: out<=0;
   49880: out<=1;
   49881: out<=1;
   49882: out<=1;
   49883: out<=1;
   49884: out<=1;
   49885: out<=0;
   49886: out<=0;
   49887: out<=1;
   49888: out<=1;
   49889: out<=0;
   49890: out<=1;
   49891: out<=0;
   49892: out<=1;
   49893: out<=1;
   49894: out<=0;
   49895: out<=0;
   49896: out<=1;
   49897: out<=1;
   49898: out<=1;
   49899: out<=1;
   49900: out<=1;
   49901: out<=0;
   49902: out<=0;
   49903: out<=1;
   49904: out<=1;
   49905: out<=0;
   49906: out<=1;
   49907: out<=0;
   49908: out<=1;
   49909: out<=1;
   49910: out<=0;
   49911: out<=0;
   49912: out<=1;
   49913: out<=1;
   49914: out<=1;
   49915: out<=1;
   49916: out<=1;
   49917: out<=0;
   49918: out<=0;
   49919: out<=1;
   49920: out<=0;
   49921: out<=0;
   49922: out<=1;
   49923: out<=1;
   49924: out<=1;
   49925: out<=0;
   49926: out<=1;
   49927: out<=0;
   49928: out<=1;
   49929: out<=0;
   49930: out<=0;
   49931: out<=1;
   49932: out<=0;
   49933: out<=0;
   49934: out<=0;
   49935: out<=0;
   49936: out<=1;
   49937: out<=1;
   49938: out<=0;
   49939: out<=0;
   49940: out<=0;
   49941: out<=1;
   49942: out<=0;
   49943: out<=1;
   49944: out<=0;
   49945: out<=1;
   49946: out<=1;
   49947: out<=0;
   49948: out<=1;
   49949: out<=1;
   49950: out<=1;
   49951: out<=1;
   49952: out<=0;
   49953: out<=0;
   49954: out<=1;
   49955: out<=1;
   49956: out<=1;
   49957: out<=0;
   49958: out<=1;
   49959: out<=0;
   49960: out<=1;
   49961: out<=0;
   49962: out<=0;
   49963: out<=1;
   49964: out<=0;
   49965: out<=0;
   49966: out<=0;
   49967: out<=0;
   49968: out<=1;
   49969: out<=1;
   49970: out<=0;
   49971: out<=0;
   49972: out<=0;
   49973: out<=1;
   49974: out<=0;
   49975: out<=1;
   49976: out<=0;
   49977: out<=1;
   49978: out<=1;
   49979: out<=0;
   49980: out<=1;
   49981: out<=1;
   49982: out<=1;
   49983: out<=1;
   49984: out<=1;
   49985: out<=1;
   49986: out<=0;
   49987: out<=0;
   49988: out<=0;
   49989: out<=1;
   49990: out<=0;
   49991: out<=1;
   49992: out<=0;
   49993: out<=1;
   49994: out<=1;
   49995: out<=0;
   49996: out<=1;
   49997: out<=1;
   49998: out<=1;
   49999: out<=1;
   50000: out<=1;
   50001: out<=1;
   50002: out<=0;
   50003: out<=0;
   50004: out<=0;
   50005: out<=1;
   50006: out<=0;
   50007: out<=1;
   50008: out<=0;
   50009: out<=1;
   50010: out<=1;
   50011: out<=0;
   50012: out<=1;
   50013: out<=1;
   50014: out<=1;
   50015: out<=1;
   50016: out<=0;
   50017: out<=0;
   50018: out<=1;
   50019: out<=1;
   50020: out<=1;
   50021: out<=0;
   50022: out<=1;
   50023: out<=0;
   50024: out<=1;
   50025: out<=0;
   50026: out<=0;
   50027: out<=1;
   50028: out<=0;
   50029: out<=0;
   50030: out<=0;
   50031: out<=0;
   50032: out<=0;
   50033: out<=0;
   50034: out<=1;
   50035: out<=1;
   50036: out<=1;
   50037: out<=0;
   50038: out<=1;
   50039: out<=0;
   50040: out<=1;
   50041: out<=0;
   50042: out<=0;
   50043: out<=1;
   50044: out<=0;
   50045: out<=0;
   50046: out<=0;
   50047: out<=0;
   50048: out<=0;
   50049: out<=0;
   50050: out<=1;
   50051: out<=1;
   50052: out<=1;
   50053: out<=0;
   50054: out<=1;
   50055: out<=0;
   50056: out<=1;
   50057: out<=0;
   50058: out<=0;
   50059: out<=1;
   50060: out<=0;
   50061: out<=0;
   50062: out<=0;
   50063: out<=0;
   50064: out<=0;
   50065: out<=0;
   50066: out<=1;
   50067: out<=1;
   50068: out<=1;
   50069: out<=0;
   50070: out<=1;
   50071: out<=0;
   50072: out<=1;
   50073: out<=0;
   50074: out<=0;
   50075: out<=1;
   50076: out<=0;
   50077: out<=0;
   50078: out<=0;
   50079: out<=0;
   50080: out<=0;
   50081: out<=0;
   50082: out<=1;
   50083: out<=1;
   50084: out<=1;
   50085: out<=0;
   50086: out<=1;
   50087: out<=0;
   50088: out<=1;
   50089: out<=0;
   50090: out<=0;
   50091: out<=1;
   50092: out<=0;
   50093: out<=0;
   50094: out<=0;
   50095: out<=0;
   50096: out<=0;
   50097: out<=0;
   50098: out<=1;
   50099: out<=1;
   50100: out<=1;
   50101: out<=0;
   50102: out<=1;
   50103: out<=0;
   50104: out<=1;
   50105: out<=0;
   50106: out<=0;
   50107: out<=1;
   50108: out<=0;
   50109: out<=0;
   50110: out<=0;
   50111: out<=0;
   50112: out<=1;
   50113: out<=1;
   50114: out<=0;
   50115: out<=0;
   50116: out<=0;
   50117: out<=1;
   50118: out<=0;
   50119: out<=1;
   50120: out<=0;
   50121: out<=1;
   50122: out<=1;
   50123: out<=0;
   50124: out<=1;
   50125: out<=1;
   50126: out<=1;
   50127: out<=1;
   50128: out<=0;
   50129: out<=0;
   50130: out<=1;
   50131: out<=1;
   50132: out<=1;
   50133: out<=0;
   50134: out<=1;
   50135: out<=0;
   50136: out<=1;
   50137: out<=0;
   50138: out<=0;
   50139: out<=1;
   50140: out<=0;
   50141: out<=0;
   50142: out<=0;
   50143: out<=0;
   50144: out<=0;
   50145: out<=0;
   50146: out<=1;
   50147: out<=1;
   50148: out<=1;
   50149: out<=0;
   50150: out<=1;
   50151: out<=0;
   50152: out<=1;
   50153: out<=0;
   50154: out<=0;
   50155: out<=1;
   50156: out<=0;
   50157: out<=0;
   50158: out<=0;
   50159: out<=0;
   50160: out<=1;
   50161: out<=1;
   50162: out<=0;
   50163: out<=0;
   50164: out<=0;
   50165: out<=1;
   50166: out<=0;
   50167: out<=1;
   50168: out<=0;
   50169: out<=1;
   50170: out<=1;
   50171: out<=0;
   50172: out<=1;
   50173: out<=1;
   50174: out<=1;
   50175: out<=1;
   50176: out<=0;
   50177: out<=1;
   50178: out<=1;
   50179: out<=0;
   50180: out<=1;
   50181: out<=1;
   50182: out<=1;
   50183: out<=1;
   50184: out<=0;
   50185: out<=0;
   50186: out<=1;
   50187: out<=1;
   50188: out<=1;
   50189: out<=0;
   50190: out<=1;
   50191: out<=0;
   50192: out<=1;
   50193: out<=0;
   50194: out<=0;
   50195: out<=1;
   50196: out<=0;
   50197: out<=0;
   50198: out<=0;
   50199: out<=0;
   50200: out<=1;
   50201: out<=1;
   50202: out<=0;
   50203: out<=0;
   50204: out<=0;
   50205: out<=1;
   50206: out<=0;
   50207: out<=1;
   50208: out<=1;
   50209: out<=0;
   50210: out<=0;
   50211: out<=1;
   50212: out<=0;
   50213: out<=0;
   50214: out<=0;
   50215: out<=0;
   50216: out<=1;
   50217: out<=1;
   50218: out<=0;
   50219: out<=0;
   50220: out<=0;
   50221: out<=1;
   50222: out<=0;
   50223: out<=1;
   50224: out<=0;
   50225: out<=1;
   50226: out<=1;
   50227: out<=0;
   50228: out<=1;
   50229: out<=1;
   50230: out<=1;
   50231: out<=1;
   50232: out<=0;
   50233: out<=0;
   50234: out<=1;
   50235: out<=1;
   50236: out<=1;
   50237: out<=0;
   50238: out<=1;
   50239: out<=0;
   50240: out<=1;
   50241: out<=0;
   50242: out<=0;
   50243: out<=1;
   50244: out<=0;
   50245: out<=0;
   50246: out<=0;
   50247: out<=0;
   50248: out<=1;
   50249: out<=1;
   50250: out<=0;
   50251: out<=0;
   50252: out<=0;
   50253: out<=1;
   50254: out<=0;
   50255: out<=1;
   50256: out<=1;
   50257: out<=0;
   50258: out<=0;
   50259: out<=1;
   50260: out<=0;
   50261: out<=0;
   50262: out<=0;
   50263: out<=0;
   50264: out<=1;
   50265: out<=1;
   50266: out<=0;
   50267: out<=0;
   50268: out<=0;
   50269: out<=1;
   50270: out<=0;
   50271: out<=1;
   50272: out<=1;
   50273: out<=0;
   50274: out<=0;
   50275: out<=1;
   50276: out<=0;
   50277: out<=0;
   50278: out<=0;
   50279: out<=0;
   50280: out<=1;
   50281: out<=1;
   50282: out<=0;
   50283: out<=0;
   50284: out<=0;
   50285: out<=1;
   50286: out<=0;
   50287: out<=1;
   50288: out<=1;
   50289: out<=0;
   50290: out<=0;
   50291: out<=1;
   50292: out<=0;
   50293: out<=0;
   50294: out<=0;
   50295: out<=0;
   50296: out<=1;
   50297: out<=1;
   50298: out<=0;
   50299: out<=0;
   50300: out<=0;
   50301: out<=1;
   50302: out<=0;
   50303: out<=1;
   50304: out<=0;
   50305: out<=1;
   50306: out<=1;
   50307: out<=0;
   50308: out<=1;
   50309: out<=1;
   50310: out<=1;
   50311: out<=1;
   50312: out<=0;
   50313: out<=0;
   50314: out<=1;
   50315: out<=1;
   50316: out<=1;
   50317: out<=0;
   50318: out<=1;
   50319: out<=0;
   50320: out<=0;
   50321: out<=1;
   50322: out<=1;
   50323: out<=0;
   50324: out<=1;
   50325: out<=1;
   50326: out<=1;
   50327: out<=1;
   50328: out<=0;
   50329: out<=0;
   50330: out<=1;
   50331: out<=1;
   50332: out<=1;
   50333: out<=0;
   50334: out<=1;
   50335: out<=0;
   50336: out<=1;
   50337: out<=0;
   50338: out<=0;
   50339: out<=1;
   50340: out<=0;
   50341: out<=0;
   50342: out<=0;
   50343: out<=0;
   50344: out<=1;
   50345: out<=1;
   50346: out<=0;
   50347: out<=0;
   50348: out<=0;
   50349: out<=1;
   50350: out<=0;
   50351: out<=1;
   50352: out<=1;
   50353: out<=0;
   50354: out<=0;
   50355: out<=1;
   50356: out<=0;
   50357: out<=0;
   50358: out<=0;
   50359: out<=0;
   50360: out<=1;
   50361: out<=1;
   50362: out<=0;
   50363: out<=0;
   50364: out<=0;
   50365: out<=1;
   50366: out<=0;
   50367: out<=1;
   50368: out<=1;
   50369: out<=0;
   50370: out<=0;
   50371: out<=1;
   50372: out<=0;
   50373: out<=0;
   50374: out<=0;
   50375: out<=0;
   50376: out<=1;
   50377: out<=1;
   50378: out<=0;
   50379: out<=0;
   50380: out<=0;
   50381: out<=1;
   50382: out<=0;
   50383: out<=1;
   50384: out<=0;
   50385: out<=1;
   50386: out<=1;
   50387: out<=0;
   50388: out<=1;
   50389: out<=1;
   50390: out<=1;
   50391: out<=1;
   50392: out<=0;
   50393: out<=0;
   50394: out<=1;
   50395: out<=1;
   50396: out<=1;
   50397: out<=0;
   50398: out<=1;
   50399: out<=0;
   50400: out<=1;
   50401: out<=0;
   50402: out<=0;
   50403: out<=1;
   50404: out<=0;
   50405: out<=0;
   50406: out<=0;
   50407: out<=0;
   50408: out<=1;
   50409: out<=1;
   50410: out<=0;
   50411: out<=0;
   50412: out<=0;
   50413: out<=1;
   50414: out<=0;
   50415: out<=1;
   50416: out<=0;
   50417: out<=1;
   50418: out<=1;
   50419: out<=0;
   50420: out<=1;
   50421: out<=1;
   50422: out<=1;
   50423: out<=1;
   50424: out<=0;
   50425: out<=0;
   50426: out<=1;
   50427: out<=1;
   50428: out<=1;
   50429: out<=0;
   50430: out<=1;
   50431: out<=0;
   50432: out<=1;
   50433: out<=1;
   50434: out<=1;
   50435: out<=1;
   50436: out<=1;
   50437: out<=0;
   50438: out<=0;
   50439: out<=1;
   50440: out<=0;
   50441: out<=1;
   50442: out<=0;
   50443: out<=1;
   50444: out<=0;
   50445: out<=0;
   50446: out<=1;
   50447: out<=1;
   50448: out<=1;
   50449: out<=1;
   50450: out<=1;
   50451: out<=1;
   50452: out<=1;
   50453: out<=0;
   50454: out<=0;
   50455: out<=1;
   50456: out<=0;
   50457: out<=1;
   50458: out<=0;
   50459: out<=1;
   50460: out<=0;
   50461: out<=0;
   50462: out<=1;
   50463: out<=1;
   50464: out<=1;
   50465: out<=1;
   50466: out<=1;
   50467: out<=1;
   50468: out<=1;
   50469: out<=0;
   50470: out<=0;
   50471: out<=1;
   50472: out<=0;
   50473: out<=1;
   50474: out<=0;
   50475: out<=1;
   50476: out<=0;
   50477: out<=0;
   50478: out<=1;
   50479: out<=1;
   50480: out<=1;
   50481: out<=1;
   50482: out<=1;
   50483: out<=1;
   50484: out<=1;
   50485: out<=0;
   50486: out<=0;
   50487: out<=1;
   50488: out<=0;
   50489: out<=1;
   50490: out<=0;
   50491: out<=1;
   50492: out<=0;
   50493: out<=0;
   50494: out<=1;
   50495: out<=1;
   50496: out<=0;
   50497: out<=0;
   50498: out<=0;
   50499: out<=0;
   50500: out<=0;
   50501: out<=1;
   50502: out<=1;
   50503: out<=0;
   50504: out<=1;
   50505: out<=0;
   50506: out<=1;
   50507: out<=0;
   50508: out<=1;
   50509: out<=1;
   50510: out<=0;
   50511: out<=0;
   50512: out<=1;
   50513: out<=1;
   50514: out<=1;
   50515: out<=1;
   50516: out<=1;
   50517: out<=0;
   50518: out<=0;
   50519: out<=1;
   50520: out<=0;
   50521: out<=1;
   50522: out<=0;
   50523: out<=1;
   50524: out<=0;
   50525: out<=0;
   50526: out<=1;
   50527: out<=1;
   50528: out<=1;
   50529: out<=1;
   50530: out<=1;
   50531: out<=1;
   50532: out<=1;
   50533: out<=0;
   50534: out<=0;
   50535: out<=1;
   50536: out<=0;
   50537: out<=1;
   50538: out<=0;
   50539: out<=1;
   50540: out<=0;
   50541: out<=0;
   50542: out<=1;
   50543: out<=1;
   50544: out<=0;
   50545: out<=0;
   50546: out<=0;
   50547: out<=0;
   50548: out<=0;
   50549: out<=1;
   50550: out<=1;
   50551: out<=0;
   50552: out<=1;
   50553: out<=0;
   50554: out<=1;
   50555: out<=0;
   50556: out<=1;
   50557: out<=1;
   50558: out<=0;
   50559: out<=0;
   50560: out<=1;
   50561: out<=1;
   50562: out<=1;
   50563: out<=1;
   50564: out<=1;
   50565: out<=0;
   50566: out<=0;
   50567: out<=1;
   50568: out<=0;
   50569: out<=1;
   50570: out<=0;
   50571: out<=1;
   50572: out<=0;
   50573: out<=0;
   50574: out<=1;
   50575: out<=1;
   50576: out<=0;
   50577: out<=0;
   50578: out<=0;
   50579: out<=0;
   50580: out<=0;
   50581: out<=1;
   50582: out<=1;
   50583: out<=0;
   50584: out<=1;
   50585: out<=0;
   50586: out<=1;
   50587: out<=0;
   50588: out<=1;
   50589: out<=1;
   50590: out<=0;
   50591: out<=0;
   50592: out<=1;
   50593: out<=1;
   50594: out<=1;
   50595: out<=1;
   50596: out<=1;
   50597: out<=0;
   50598: out<=0;
   50599: out<=1;
   50600: out<=0;
   50601: out<=1;
   50602: out<=0;
   50603: out<=1;
   50604: out<=0;
   50605: out<=0;
   50606: out<=1;
   50607: out<=1;
   50608: out<=0;
   50609: out<=0;
   50610: out<=0;
   50611: out<=0;
   50612: out<=0;
   50613: out<=1;
   50614: out<=1;
   50615: out<=0;
   50616: out<=1;
   50617: out<=0;
   50618: out<=1;
   50619: out<=0;
   50620: out<=1;
   50621: out<=1;
   50622: out<=0;
   50623: out<=0;
   50624: out<=0;
   50625: out<=0;
   50626: out<=0;
   50627: out<=0;
   50628: out<=0;
   50629: out<=1;
   50630: out<=1;
   50631: out<=0;
   50632: out<=1;
   50633: out<=0;
   50634: out<=1;
   50635: out<=0;
   50636: out<=1;
   50637: out<=1;
   50638: out<=0;
   50639: out<=0;
   50640: out<=0;
   50641: out<=0;
   50642: out<=0;
   50643: out<=0;
   50644: out<=0;
   50645: out<=1;
   50646: out<=1;
   50647: out<=0;
   50648: out<=1;
   50649: out<=0;
   50650: out<=1;
   50651: out<=0;
   50652: out<=1;
   50653: out<=1;
   50654: out<=0;
   50655: out<=0;
   50656: out<=1;
   50657: out<=1;
   50658: out<=1;
   50659: out<=1;
   50660: out<=1;
   50661: out<=0;
   50662: out<=0;
   50663: out<=1;
   50664: out<=0;
   50665: out<=1;
   50666: out<=0;
   50667: out<=1;
   50668: out<=0;
   50669: out<=0;
   50670: out<=1;
   50671: out<=1;
   50672: out<=1;
   50673: out<=1;
   50674: out<=1;
   50675: out<=1;
   50676: out<=1;
   50677: out<=0;
   50678: out<=0;
   50679: out<=1;
   50680: out<=0;
   50681: out<=1;
   50682: out<=0;
   50683: out<=1;
   50684: out<=0;
   50685: out<=0;
   50686: out<=1;
   50687: out<=1;
   50688: out<=1;
   50689: out<=1;
   50690: out<=0;
   50691: out<=0;
   50692: out<=1;
   50693: out<=0;
   50694: out<=1;
   50695: out<=0;
   50696: out<=1;
   50697: out<=0;
   50698: out<=0;
   50699: out<=1;
   50700: out<=1;
   50701: out<=1;
   50702: out<=1;
   50703: out<=1;
   50704: out<=1;
   50705: out<=1;
   50706: out<=0;
   50707: out<=0;
   50708: out<=1;
   50709: out<=0;
   50710: out<=1;
   50711: out<=0;
   50712: out<=1;
   50713: out<=0;
   50714: out<=0;
   50715: out<=1;
   50716: out<=1;
   50717: out<=1;
   50718: out<=1;
   50719: out<=1;
   50720: out<=0;
   50721: out<=0;
   50722: out<=1;
   50723: out<=1;
   50724: out<=0;
   50725: out<=1;
   50726: out<=0;
   50727: out<=1;
   50728: out<=0;
   50729: out<=1;
   50730: out<=1;
   50731: out<=0;
   50732: out<=0;
   50733: out<=0;
   50734: out<=0;
   50735: out<=0;
   50736: out<=0;
   50737: out<=0;
   50738: out<=1;
   50739: out<=1;
   50740: out<=0;
   50741: out<=1;
   50742: out<=0;
   50743: out<=1;
   50744: out<=0;
   50745: out<=1;
   50746: out<=1;
   50747: out<=0;
   50748: out<=0;
   50749: out<=0;
   50750: out<=0;
   50751: out<=0;
   50752: out<=0;
   50753: out<=0;
   50754: out<=1;
   50755: out<=1;
   50756: out<=0;
   50757: out<=1;
   50758: out<=0;
   50759: out<=1;
   50760: out<=0;
   50761: out<=1;
   50762: out<=1;
   50763: out<=0;
   50764: out<=0;
   50765: out<=0;
   50766: out<=0;
   50767: out<=0;
   50768: out<=1;
   50769: out<=1;
   50770: out<=0;
   50771: out<=0;
   50772: out<=1;
   50773: out<=0;
   50774: out<=1;
   50775: out<=0;
   50776: out<=1;
   50777: out<=0;
   50778: out<=0;
   50779: out<=1;
   50780: out<=1;
   50781: out<=1;
   50782: out<=1;
   50783: out<=1;
   50784: out<=0;
   50785: out<=0;
   50786: out<=1;
   50787: out<=1;
   50788: out<=0;
   50789: out<=1;
   50790: out<=0;
   50791: out<=1;
   50792: out<=0;
   50793: out<=1;
   50794: out<=1;
   50795: out<=0;
   50796: out<=0;
   50797: out<=0;
   50798: out<=0;
   50799: out<=0;
   50800: out<=1;
   50801: out<=1;
   50802: out<=0;
   50803: out<=0;
   50804: out<=1;
   50805: out<=0;
   50806: out<=1;
   50807: out<=0;
   50808: out<=1;
   50809: out<=0;
   50810: out<=0;
   50811: out<=1;
   50812: out<=1;
   50813: out<=1;
   50814: out<=1;
   50815: out<=1;
   50816: out<=1;
   50817: out<=1;
   50818: out<=0;
   50819: out<=0;
   50820: out<=1;
   50821: out<=0;
   50822: out<=1;
   50823: out<=0;
   50824: out<=1;
   50825: out<=0;
   50826: out<=0;
   50827: out<=1;
   50828: out<=1;
   50829: out<=1;
   50830: out<=1;
   50831: out<=1;
   50832: out<=0;
   50833: out<=0;
   50834: out<=1;
   50835: out<=1;
   50836: out<=0;
   50837: out<=1;
   50838: out<=0;
   50839: out<=1;
   50840: out<=0;
   50841: out<=1;
   50842: out<=1;
   50843: out<=0;
   50844: out<=0;
   50845: out<=0;
   50846: out<=0;
   50847: out<=0;
   50848: out<=0;
   50849: out<=0;
   50850: out<=1;
   50851: out<=1;
   50852: out<=0;
   50853: out<=1;
   50854: out<=0;
   50855: out<=1;
   50856: out<=0;
   50857: out<=1;
   50858: out<=1;
   50859: out<=0;
   50860: out<=0;
   50861: out<=0;
   50862: out<=0;
   50863: out<=0;
   50864: out<=1;
   50865: out<=1;
   50866: out<=0;
   50867: out<=0;
   50868: out<=1;
   50869: out<=0;
   50870: out<=1;
   50871: out<=0;
   50872: out<=1;
   50873: out<=0;
   50874: out<=0;
   50875: out<=1;
   50876: out<=1;
   50877: out<=1;
   50878: out<=1;
   50879: out<=1;
   50880: out<=0;
   50881: out<=0;
   50882: out<=1;
   50883: out<=1;
   50884: out<=0;
   50885: out<=1;
   50886: out<=0;
   50887: out<=1;
   50888: out<=0;
   50889: out<=1;
   50890: out<=1;
   50891: out<=0;
   50892: out<=0;
   50893: out<=0;
   50894: out<=0;
   50895: out<=0;
   50896: out<=0;
   50897: out<=0;
   50898: out<=1;
   50899: out<=1;
   50900: out<=0;
   50901: out<=1;
   50902: out<=0;
   50903: out<=1;
   50904: out<=0;
   50905: out<=1;
   50906: out<=1;
   50907: out<=0;
   50908: out<=0;
   50909: out<=0;
   50910: out<=0;
   50911: out<=0;
   50912: out<=0;
   50913: out<=0;
   50914: out<=1;
   50915: out<=1;
   50916: out<=0;
   50917: out<=1;
   50918: out<=0;
   50919: out<=1;
   50920: out<=0;
   50921: out<=1;
   50922: out<=1;
   50923: out<=0;
   50924: out<=0;
   50925: out<=0;
   50926: out<=0;
   50927: out<=0;
   50928: out<=0;
   50929: out<=0;
   50930: out<=1;
   50931: out<=1;
   50932: out<=0;
   50933: out<=1;
   50934: out<=0;
   50935: out<=1;
   50936: out<=0;
   50937: out<=1;
   50938: out<=1;
   50939: out<=0;
   50940: out<=0;
   50941: out<=0;
   50942: out<=0;
   50943: out<=0;
   50944: out<=0;
   50945: out<=1;
   50946: out<=0;
   50947: out<=1;
   50948: out<=1;
   50949: out<=1;
   50950: out<=0;
   50951: out<=0;
   50952: out<=1;
   50953: out<=1;
   50954: out<=1;
   50955: out<=1;
   50956: out<=0;
   50957: out<=1;
   50958: out<=1;
   50959: out<=0;
   50960: out<=1;
   50961: out<=0;
   50962: out<=1;
   50963: out<=0;
   50964: out<=0;
   50965: out<=0;
   50966: out<=1;
   50967: out<=1;
   50968: out<=0;
   50969: out<=0;
   50970: out<=0;
   50971: out<=0;
   50972: out<=1;
   50973: out<=0;
   50974: out<=0;
   50975: out<=1;
   50976: out<=0;
   50977: out<=1;
   50978: out<=0;
   50979: out<=1;
   50980: out<=1;
   50981: out<=1;
   50982: out<=0;
   50983: out<=0;
   50984: out<=1;
   50985: out<=1;
   50986: out<=1;
   50987: out<=1;
   50988: out<=0;
   50989: out<=1;
   50990: out<=1;
   50991: out<=0;
   50992: out<=1;
   50993: out<=0;
   50994: out<=1;
   50995: out<=0;
   50996: out<=0;
   50997: out<=0;
   50998: out<=1;
   50999: out<=1;
   51000: out<=0;
   51001: out<=0;
   51002: out<=0;
   51003: out<=0;
   51004: out<=1;
   51005: out<=0;
   51006: out<=0;
   51007: out<=1;
   51008: out<=1;
   51009: out<=0;
   51010: out<=1;
   51011: out<=0;
   51012: out<=0;
   51013: out<=0;
   51014: out<=1;
   51015: out<=1;
   51016: out<=0;
   51017: out<=0;
   51018: out<=0;
   51019: out<=0;
   51020: out<=1;
   51021: out<=0;
   51022: out<=0;
   51023: out<=1;
   51024: out<=1;
   51025: out<=0;
   51026: out<=1;
   51027: out<=0;
   51028: out<=0;
   51029: out<=0;
   51030: out<=1;
   51031: out<=1;
   51032: out<=0;
   51033: out<=0;
   51034: out<=0;
   51035: out<=0;
   51036: out<=1;
   51037: out<=0;
   51038: out<=0;
   51039: out<=1;
   51040: out<=0;
   51041: out<=1;
   51042: out<=0;
   51043: out<=1;
   51044: out<=1;
   51045: out<=1;
   51046: out<=0;
   51047: out<=0;
   51048: out<=1;
   51049: out<=1;
   51050: out<=1;
   51051: out<=1;
   51052: out<=0;
   51053: out<=1;
   51054: out<=1;
   51055: out<=0;
   51056: out<=0;
   51057: out<=1;
   51058: out<=0;
   51059: out<=1;
   51060: out<=1;
   51061: out<=1;
   51062: out<=0;
   51063: out<=0;
   51064: out<=1;
   51065: out<=1;
   51066: out<=1;
   51067: out<=1;
   51068: out<=0;
   51069: out<=1;
   51070: out<=1;
   51071: out<=0;
   51072: out<=0;
   51073: out<=1;
   51074: out<=0;
   51075: out<=1;
   51076: out<=1;
   51077: out<=1;
   51078: out<=0;
   51079: out<=0;
   51080: out<=1;
   51081: out<=1;
   51082: out<=1;
   51083: out<=1;
   51084: out<=0;
   51085: out<=1;
   51086: out<=1;
   51087: out<=0;
   51088: out<=0;
   51089: out<=1;
   51090: out<=0;
   51091: out<=1;
   51092: out<=1;
   51093: out<=1;
   51094: out<=0;
   51095: out<=0;
   51096: out<=1;
   51097: out<=1;
   51098: out<=1;
   51099: out<=1;
   51100: out<=0;
   51101: out<=1;
   51102: out<=1;
   51103: out<=0;
   51104: out<=0;
   51105: out<=1;
   51106: out<=0;
   51107: out<=1;
   51108: out<=1;
   51109: out<=1;
   51110: out<=0;
   51111: out<=0;
   51112: out<=1;
   51113: out<=1;
   51114: out<=1;
   51115: out<=1;
   51116: out<=0;
   51117: out<=1;
   51118: out<=1;
   51119: out<=0;
   51120: out<=0;
   51121: out<=1;
   51122: out<=0;
   51123: out<=1;
   51124: out<=1;
   51125: out<=1;
   51126: out<=0;
   51127: out<=0;
   51128: out<=1;
   51129: out<=1;
   51130: out<=1;
   51131: out<=1;
   51132: out<=0;
   51133: out<=1;
   51134: out<=1;
   51135: out<=0;
   51136: out<=1;
   51137: out<=0;
   51138: out<=1;
   51139: out<=0;
   51140: out<=0;
   51141: out<=0;
   51142: out<=1;
   51143: out<=1;
   51144: out<=0;
   51145: out<=0;
   51146: out<=0;
   51147: out<=0;
   51148: out<=1;
   51149: out<=0;
   51150: out<=0;
   51151: out<=1;
   51152: out<=0;
   51153: out<=1;
   51154: out<=0;
   51155: out<=1;
   51156: out<=1;
   51157: out<=1;
   51158: out<=0;
   51159: out<=0;
   51160: out<=1;
   51161: out<=1;
   51162: out<=1;
   51163: out<=1;
   51164: out<=0;
   51165: out<=1;
   51166: out<=1;
   51167: out<=0;
   51168: out<=0;
   51169: out<=1;
   51170: out<=0;
   51171: out<=1;
   51172: out<=1;
   51173: out<=1;
   51174: out<=0;
   51175: out<=0;
   51176: out<=1;
   51177: out<=1;
   51178: out<=1;
   51179: out<=1;
   51180: out<=0;
   51181: out<=1;
   51182: out<=1;
   51183: out<=0;
   51184: out<=1;
   51185: out<=0;
   51186: out<=1;
   51187: out<=0;
   51188: out<=0;
   51189: out<=0;
   51190: out<=1;
   51191: out<=1;
   51192: out<=0;
   51193: out<=0;
   51194: out<=0;
   51195: out<=0;
   51196: out<=1;
   51197: out<=0;
   51198: out<=0;
   51199: out<=1;
   51200: out<=0;
   51201: out<=1;
   51202: out<=0;
   51203: out<=1;
   51204: out<=1;
   51205: out<=1;
   51206: out<=0;
   51207: out<=0;
   51208: out<=0;
   51209: out<=0;
   51210: out<=0;
   51211: out<=0;
   51212: out<=1;
   51213: out<=0;
   51214: out<=0;
   51215: out<=1;
   51216: out<=1;
   51217: out<=0;
   51218: out<=1;
   51219: out<=0;
   51220: out<=0;
   51221: out<=0;
   51222: out<=1;
   51223: out<=1;
   51224: out<=1;
   51225: out<=1;
   51226: out<=1;
   51227: out<=1;
   51228: out<=0;
   51229: out<=1;
   51230: out<=1;
   51231: out<=0;
   51232: out<=1;
   51233: out<=0;
   51234: out<=1;
   51235: out<=0;
   51236: out<=0;
   51237: out<=0;
   51238: out<=1;
   51239: out<=1;
   51240: out<=1;
   51241: out<=1;
   51242: out<=1;
   51243: out<=1;
   51244: out<=0;
   51245: out<=1;
   51246: out<=1;
   51247: out<=0;
   51248: out<=0;
   51249: out<=1;
   51250: out<=0;
   51251: out<=1;
   51252: out<=1;
   51253: out<=1;
   51254: out<=0;
   51255: out<=0;
   51256: out<=0;
   51257: out<=0;
   51258: out<=0;
   51259: out<=0;
   51260: out<=1;
   51261: out<=0;
   51262: out<=0;
   51263: out<=1;
   51264: out<=1;
   51265: out<=0;
   51266: out<=1;
   51267: out<=0;
   51268: out<=0;
   51269: out<=0;
   51270: out<=1;
   51271: out<=1;
   51272: out<=1;
   51273: out<=1;
   51274: out<=1;
   51275: out<=1;
   51276: out<=0;
   51277: out<=1;
   51278: out<=1;
   51279: out<=0;
   51280: out<=1;
   51281: out<=0;
   51282: out<=1;
   51283: out<=0;
   51284: out<=0;
   51285: out<=0;
   51286: out<=1;
   51287: out<=1;
   51288: out<=1;
   51289: out<=1;
   51290: out<=1;
   51291: out<=1;
   51292: out<=0;
   51293: out<=1;
   51294: out<=1;
   51295: out<=0;
   51296: out<=1;
   51297: out<=0;
   51298: out<=1;
   51299: out<=0;
   51300: out<=0;
   51301: out<=0;
   51302: out<=1;
   51303: out<=1;
   51304: out<=1;
   51305: out<=1;
   51306: out<=1;
   51307: out<=1;
   51308: out<=0;
   51309: out<=1;
   51310: out<=1;
   51311: out<=0;
   51312: out<=1;
   51313: out<=0;
   51314: out<=1;
   51315: out<=0;
   51316: out<=0;
   51317: out<=0;
   51318: out<=1;
   51319: out<=1;
   51320: out<=1;
   51321: out<=1;
   51322: out<=1;
   51323: out<=1;
   51324: out<=0;
   51325: out<=1;
   51326: out<=1;
   51327: out<=0;
   51328: out<=0;
   51329: out<=1;
   51330: out<=0;
   51331: out<=1;
   51332: out<=1;
   51333: out<=1;
   51334: out<=0;
   51335: out<=0;
   51336: out<=0;
   51337: out<=0;
   51338: out<=0;
   51339: out<=0;
   51340: out<=1;
   51341: out<=0;
   51342: out<=0;
   51343: out<=1;
   51344: out<=0;
   51345: out<=1;
   51346: out<=0;
   51347: out<=1;
   51348: out<=1;
   51349: out<=1;
   51350: out<=0;
   51351: out<=0;
   51352: out<=0;
   51353: out<=0;
   51354: out<=0;
   51355: out<=0;
   51356: out<=1;
   51357: out<=0;
   51358: out<=0;
   51359: out<=1;
   51360: out<=1;
   51361: out<=0;
   51362: out<=1;
   51363: out<=0;
   51364: out<=0;
   51365: out<=0;
   51366: out<=1;
   51367: out<=1;
   51368: out<=1;
   51369: out<=1;
   51370: out<=1;
   51371: out<=1;
   51372: out<=0;
   51373: out<=1;
   51374: out<=1;
   51375: out<=0;
   51376: out<=1;
   51377: out<=0;
   51378: out<=1;
   51379: out<=0;
   51380: out<=0;
   51381: out<=0;
   51382: out<=1;
   51383: out<=1;
   51384: out<=1;
   51385: out<=1;
   51386: out<=1;
   51387: out<=1;
   51388: out<=0;
   51389: out<=1;
   51390: out<=1;
   51391: out<=0;
   51392: out<=1;
   51393: out<=0;
   51394: out<=1;
   51395: out<=0;
   51396: out<=0;
   51397: out<=0;
   51398: out<=1;
   51399: out<=1;
   51400: out<=1;
   51401: out<=1;
   51402: out<=1;
   51403: out<=1;
   51404: out<=0;
   51405: out<=1;
   51406: out<=1;
   51407: out<=0;
   51408: out<=0;
   51409: out<=1;
   51410: out<=0;
   51411: out<=1;
   51412: out<=1;
   51413: out<=1;
   51414: out<=0;
   51415: out<=0;
   51416: out<=0;
   51417: out<=0;
   51418: out<=0;
   51419: out<=0;
   51420: out<=1;
   51421: out<=0;
   51422: out<=0;
   51423: out<=1;
   51424: out<=1;
   51425: out<=0;
   51426: out<=1;
   51427: out<=0;
   51428: out<=0;
   51429: out<=0;
   51430: out<=1;
   51431: out<=1;
   51432: out<=1;
   51433: out<=1;
   51434: out<=1;
   51435: out<=1;
   51436: out<=0;
   51437: out<=1;
   51438: out<=1;
   51439: out<=0;
   51440: out<=0;
   51441: out<=1;
   51442: out<=0;
   51443: out<=1;
   51444: out<=1;
   51445: out<=1;
   51446: out<=0;
   51447: out<=0;
   51448: out<=0;
   51449: out<=0;
   51450: out<=0;
   51451: out<=0;
   51452: out<=1;
   51453: out<=0;
   51454: out<=0;
   51455: out<=1;
   51456: out<=1;
   51457: out<=1;
   51458: out<=0;
   51459: out<=0;
   51460: out<=1;
   51461: out<=0;
   51462: out<=1;
   51463: out<=0;
   51464: out<=0;
   51465: out<=1;
   51466: out<=1;
   51467: out<=0;
   51468: out<=0;
   51469: out<=0;
   51470: out<=0;
   51471: out<=0;
   51472: out<=1;
   51473: out<=1;
   51474: out<=0;
   51475: out<=0;
   51476: out<=1;
   51477: out<=0;
   51478: out<=1;
   51479: out<=0;
   51480: out<=0;
   51481: out<=1;
   51482: out<=1;
   51483: out<=0;
   51484: out<=0;
   51485: out<=0;
   51486: out<=0;
   51487: out<=0;
   51488: out<=1;
   51489: out<=1;
   51490: out<=0;
   51491: out<=0;
   51492: out<=1;
   51493: out<=0;
   51494: out<=1;
   51495: out<=0;
   51496: out<=0;
   51497: out<=1;
   51498: out<=1;
   51499: out<=0;
   51500: out<=0;
   51501: out<=0;
   51502: out<=0;
   51503: out<=0;
   51504: out<=1;
   51505: out<=1;
   51506: out<=0;
   51507: out<=0;
   51508: out<=1;
   51509: out<=0;
   51510: out<=1;
   51511: out<=0;
   51512: out<=0;
   51513: out<=1;
   51514: out<=1;
   51515: out<=0;
   51516: out<=0;
   51517: out<=0;
   51518: out<=0;
   51519: out<=0;
   51520: out<=0;
   51521: out<=0;
   51522: out<=1;
   51523: out<=1;
   51524: out<=0;
   51525: out<=1;
   51526: out<=0;
   51527: out<=1;
   51528: out<=1;
   51529: out<=0;
   51530: out<=0;
   51531: out<=1;
   51532: out<=1;
   51533: out<=1;
   51534: out<=1;
   51535: out<=1;
   51536: out<=1;
   51537: out<=1;
   51538: out<=0;
   51539: out<=0;
   51540: out<=1;
   51541: out<=0;
   51542: out<=1;
   51543: out<=0;
   51544: out<=0;
   51545: out<=1;
   51546: out<=1;
   51547: out<=0;
   51548: out<=0;
   51549: out<=0;
   51550: out<=0;
   51551: out<=0;
   51552: out<=1;
   51553: out<=1;
   51554: out<=0;
   51555: out<=0;
   51556: out<=1;
   51557: out<=0;
   51558: out<=1;
   51559: out<=0;
   51560: out<=0;
   51561: out<=1;
   51562: out<=1;
   51563: out<=0;
   51564: out<=0;
   51565: out<=0;
   51566: out<=0;
   51567: out<=0;
   51568: out<=0;
   51569: out<=0;
   51570: out<=1;
   51571: out<=1;
   51572: out<=0;
   51573: out<=1;
   51574: out<=0;
   51575: out<=1;
   51576: out<=1;
   51577: out<=0;
   51578: out<=0;
   51579: out<=1;
   51580: out<=1;
   51581: out<=1;
   51582: out<=1;
   51583: out<=1;
   51584: out<=1;
   51585: out<=1;
   51586: out<=0;
   51587: out<=0;
   51588: out<=1;
   51589: out<=0;
   51590: out<=1;
   51591: out<=0;
   51592: out<=0;
   51593: out<=1;
   51594: out<=1;
   51595: out<=0;
   51596: out<=0;
   51597: out<=0;
   51598: out<=0;
   51599: out<=0;
   51600: out<=0;
   51601: out<=0;
   51602: out<=1;
   51603: out<=1;
   51604: out<=0;
   51605: out<=1;
   51606: out<=0;
   51607: out<=1;
   51608: out<=1;
   51609: out<=0;
   51610: out<=0;
   51611: out<=1;
   51612: out<=1;
   51613: out<=1;
   51614: out<=1;
   51615: out<=1;
   51616: out<=1;
   51617: out<=1;
   51618: out<=0;
   51619: out<=0;
   51620: out<=1;
   51621: out<=0;
   51622: out<=1;
   51623: out<=0;
   51624: out<=0;
   51625: out<=1;
   51626: out<=1;
   51627: out<=0;
   51628: out<=0;
   51629: out<=0;
   51630: out<=0;
   51631: out<=0;
   51632: out<=0;
   51633: out<=0;
   51634: out<=1;
   51635: out<=1;
   51636: out<=0;
   51637: out<=1;
   51638: out<=0;
   51639: out<=1;
   51640: out<=1;
   51641: out<=0;
   51642: out<=0;
   51643: out<=1;
   51644: out<=1;
   51645: out<=1;
   51646: out<=1;
   51647: out<=1;
   51648: out<=0;
   51649: out<=0;
   51650: out<=1;
   51651: out<=1;
   51652: out<=0;
   51653: out<=1;
   51654: out<=0;
   51655: out<=1;
   51656: out<=1;
   51657: out<=0;
   51658: out<=0;
   51659: out<=1;
   51660: out<=1;
   51661: out<=1;
   51662: out<=1;
   51663: out<=1;
   51664: out<=0;
   51665: out<=0;
   51666: out<=1;
   51667: out<=1;
   51668: out<=0;
   51669: out<=1;
   51670: out<=0;
   51671: out<=1;
   51672: out<=1;
   51673: out<=0;
   51674: out<=0;
   51675: out<=1;
   51676: out<=1;
   51677: out<=1;
   51678: out<=1;
   51679: out<=1;
   51680: out<=1;
   51681: out<=1;
   51682: out<=0;
   51683: out<=0;
   51684: out<=1;
   51685: out<=0;
   51686: out<=1;
   51687: out<=0;
   51688: out<=0;
   51689: out<=1;
   51690: out<=1;
   51691: out<=0;
   51692: out<=0;
   51693: out<=0;
   51694: out<=0;
   51695: out<=0;
   51696: out<=1;
   51697: out<=1;
   51698: out<=0;
   51699: out<=0;
   51700: out<=1;
   51701: out<=0;
   51702: out<=1;
   51703: out<=0;
   51704: out<=0;
   51705: out<=1;
   51706: out<=1;
   51707: out<=0;
   51708: out<=0;
   51709: out<=0;
   51710: out<=0;
   51711: out<=0;
   51712: out<=0;
   51713: out<=0;
   51714: out<=0;
   51715: out<=0;
   51716: out<=0;
   51717: out<=1;
   51718: out<=1;
   51719: out<=0;
   51720: out<=0;
   51721: out<=1;
   51722: out<=0;
   51723: out<=1;
   51724: out<=0;
   51725: out<=0;
   51726: out<=1;
   51727: out<=1;
   51728: out<=0;
   51729: out<=0;
   51730: out<=0;
   51731: out<=0;
   51732: out<=0;
   51733: out<=1;
   51734: out<=1;
   51735: out<=0;
   51736: out<=0;
   51737: out<=1;
   51738: out<=0;
   51739: out<=1;
   51740: out<=0;
   51741: out<=0;
   51742: out<=1;
   51743: out<=1;
   51744: out<=1;
   51745: out<=1;
   51746: out<=1;
   51747: out<=1;
   51748: out<=1;
   51749: out<=0;
   51750: out<=0;
   51751: out<=1;
   51752: out<=1;
   51753: out<=0;
   51754: out<=1;
   51755: out<=0;
   51756: out<=1;
   51757: out<=1;
   51758: out<=0;
   51759: out<=0;
   51760: out<=1;
   51761: out<=1;
   51762: out<=1;
   51763: out<=1;
   51764: out<=1;
   51765: out<=0;
   51766: out<=0;
   51767: out<=1;
   51768: out<=1;
   51769: out<=0;
   51770: out<=1;
   51771: out<=0;
   51772: out<=1;
   51773: out<=1;
   51774: out<=0;
   51775: out<=0;
   51776: out<=1;
   51777: out<=1;
   51778: out<=1;
   51779: out<=1;
   51780: out<=1;
   51781: out<=0;
   51782: out<=0;
   51783: out<=1;
   51784: out<=1;
   51785: out<=0;
   51786: out<=1;
   51787: out<=0;
   51788: out<=1;
   51789: out<=1;
   51790: out<=0;
   51791: out<=0;
   51792: out<=0;
   51793: out<=0;
   51794: out<=0;
   51795: out<=0;
   51796: out<=0;
   51797: out<=1;
   51798: out<=1;
   51799: out<=0;
   51800: out<=0;
   51801: out<=1;
   51802: out<=0;
   51803: out<=1;
   51804: out<=0;
   51805: out<=0;
   51806: out<=1;
   51807: out<=1;
   51808: out<=1;
   51809: out<=1;
   51810: out<=1;
   51811: out<=1;
   51812: out<=1;
   51813: out<=0;
   51814: out<=0;
   51815: out<=1;
   51816: out<=1;
   51817: out<=0;
   51818: out<=1;
   51819: out<=0;
   51820: out<=1;
   51821: out<=1;
   51822: out<=0;
   51823: out<=0;
   51824: out<=0;
   51825: out<=0;
   51826: out<=0;
   51827: out<=0;
   51828: out<=0;
   51829: out<=1;
   51830: out<=1;
   51831: out<=0;
   51832: out<=0;
   51833: out<=1;
   51834: out<=0;
   51835: out<=1;
   51836: out<=0;
   51837: out<=0;
   51838: out<=1;
   51839: out<=1;
   51840: out<=0;
   51841: out<=0;
   51842: out<=0;
   51843: out<=0;
   51844: out<=0;
   51845: out<=1;
   51846: out<=1;
   51847: out<=0;
   51848: out<=0;
   51849: out<=1;
   51850: out<=0;
   51851: out<=1;
   51852: out<=0;
   51853: out<=0;
   51854: out<=1;
   51855: out<=1;
   51856: out<=1;
   51857: out<=1;
   51858: out<=1;
   51859: out<=1;
   51860: out<=1;
   51861: out<=0;
   51862: out<=0;
   51863: out<=1;
   51864: out<=1;
   51865: out<=0;
   51866: out<=1;
   51867: out<=0;
   51868: out<=1;
   51869: out<=1;
   51870: out<=0;
   51871: out<=0;
   51872: out<=1;
   51873: out<=1;
   51874: out<=1;
   51875: out<=1;
   51876: out<=1;
   51877: out<=0;
   51878: out<=0;
   51879: out<=1;
   51880: out<=1;
   51881: out<=0;
   51882: out<=1;
   51883: out<=0;
   51884: out<=1;
   51885: out<=1;
   51886: out<=0;
   51887: out<=0;
   51888: out<=0;
   51889: out<=0;
   51890: out<=0;
   51891: out<=0;
   51892: out<=0;
   51893: out<=1;
   51894: out<=1;
   51895: out<=0;
   51896: out<=0;
   51897: out<=1;
   51898: out<=0;
   51899: out<=1;
   51900: out<=0;
   51901: out<=0;
   51902: out<=1;
   51903: out<=1;
   51904: out<=1;
   51905: out<=1;
   51906: out<=1;
   51907: out<=1;
   51908: out<=1;
   51909: out<=0;
   51910: out<=0;
   51911: out<=1;
   51912: out<=1;
   51913: out<=0;
   51914: out<=1;
   51915: out<=0;
   51916: out<=1;
   51917: out<=1;
   51918: out<=0;
   51919: out<=0;
   51920: out<=1;
   51921: out<=1;
   51922: out<=1;
   51923: out<=1;
   51924: out<=1;
   51925: out<=0;
   51926: out<=0;
   51927: out<=1;
   51928: out<=1;
   51929: out<=0;
   51930: out<=1;
   51931: out<=0;
   51932: out<=1;
   51933: out<=1;
   51934: out<=0;
   51935: out<=0;
   51936: out<=1;
   51937: out<=1;
   51938: out<=1;
   51939: out<=1;
   51940: out<=1;
   51941: out<=0;
   51942: out<=0;
   51943: out<=1;
   51944: out<=1;
   51945: out<=0;
   51946: out<=1;
   51947: out<=0;
   51948: out<=1;
   51949: out<=1;
   51950: out<=0;
   51951: out<=0;
   51952: out<=1;
   51953: out<=1;
   51954: out<=1;
   51955: out<=1;
   51956: out<=1;
   51957: out<=0;
   51958: out<=0;
   51959: out<=1;
   51960: out<=1;
   51961: out<=0;
   51962: out<=1;
   51963: out<=0;
   51964: out<=1;
   51965: out<=1;
   51966: out<=0;
   51967: out<=0;
   51968: out<=1;
   51969: out<=0;
   51970: out<=0;
   51971: out<=1;
   51972: out<=0;
   51973: out<=0;
   51974: out<=0;
   51975: out<=0;
   51976: out<=0;
   51977: out<=0;
   51978: out<=1;
   51979: out<=1;
   51980: out<=1;
   51981: out<=0;
   51982: out<=1;
   51983: out<=0;
   51984: out<=0;
   51985: out<=1;
   51986: out<=1;
   51987: out<=0;
   51988: out<=1;
   51989: out<=1;
   51990: out<=1;
   51991: out<=1;
   51992: out<=1;
   51993: out<=1;
   51994: out<=0;
   51995: out<=0;
   51996: out<=0;
   51997: out<=1;
   51998: out<=0;
   51999: out<=1;
   52000: out<=1;
   52001: out<=0;
   52002: out<=0;
   52003: out<=1;
   52004: out<=0;
   52005: out<=0;
   52006: out<=0;
   52007: out<=0;
   52008: out<=0;
   52009: out<=0;
   52010: out<=1;
   52011: out<=1;
   52012: out<=1;
   52013: out<=0;
   52014: out<=1;
   52015: out<=0;
   52016: out<=0;
   52017: out<=1;
   52018: out<=1;
   52019: out<=0;
   52020: out<=1;
   52021: out<=1;
   52022: out<=1;
   52023: out<=1;
   52024: out<=1;
   52025: out<=1;
   52026: out<=0;
   52027: out<=0;
   52028: out<=0;
   52029: out<=1;
   52030: out<=0;
   52031: out<=1;
   52032: out<=0;
   52033: out<=1;
   52034: out<=1;
   52035: out<=0;
   52036: out<=1;
   52037: out<=1;
   52038: out<=1;
   52039: out<=1;
   52040: out<=1;
   52041: out<=1;
   52042: out<=0;
   52043: out<=0;
   52044: out<=0;
   52045: out<=1;
   52046: out<=0;
   52047: out<=1;
   52048: out<=0;
   52049: out<=1;
   52050: out<=1;
   52051: out<=0;
   52052: out<=1;
   52053: out<=1;
   52054: out<=1;
   52055: out<=1;
   52056: out<=1;
   52057: out<=1;
   52058: out<=0;
   52059: out<=0;
   52060: out<=0;
   52061: out<=1;
   52062: out<=0;
   52063: out<=1;
   52064: out<=1;
   52065: out<=0;
   52066: out<=0;
   52067: out<=1;
   52068: out<=0;
   52069: out<=0;
   52070: out<=0;
   52071: out<=0;
   52072: out<=0;
   52073: out<=0;
   52074: out<=1;
   52075: out<=1;
   52076: out<=1;
   52077: out<=0;
   52078: out<=1;
   52079: out<=0;
   52080: out<=1;
   52081: out<=0;
   52082: out<=0;
   52083: out<=1;
   52084: out<=0;
   52085: out<=0;
   52086: out<=0;
   52087: out<=0;
   52088: out<=0;
   52089: out<=0;
   52090: out<=1;
   52091: out<=1;
   52092: out<=1;
   52093: out<=0;
   52094: out<=1;
   52095: out<=0;
   52096: out<=1;
   52097: out<=0;
   52098: out<=0;
   52099: out<=1;
   52100: out<=0;
   52101: out<=0;
   52102: out<=0;
   52103: out<=0;
   52104: out<=0;
   52105: out<=0;
   52106: out<=1;
   52107: out<=1;
   52108: out<=1;
   52109: out<=0;
   52110: out<=1;
   52111: out<=0;
   52112: out<=1;
   52113: out<=0;
   52114: out<=0;
   52115: out<=1;
   52116: out<=0;
   52117: out<=0;
   52118: out<=0;
   52119: out<=0;
   52120: out<=0;
   52121: out<=0;
   52122: out<=1;
   52123: out<=1;
   52124: out<=1;
   52125: out<=0;
   52126: out<=1;
   52127: out<=0;
   52128: out<=1;
   52129: out<=0;
   52130: out<=0;
   52131: out<=1;
   52132: out<=0;
   52133: out<=0;
   52134: out<=0;
   52135: out<=0;
   52136: out<=0;
   52137: out<=0;
   52138: out<=1;
   52139: out<=1;
   52140: out<=1;
   52141: out<=0;
   52142: out<=1;
   52143: out<=0;
   52144: out<=1;
   52145: out<=0;
   52146: out<=0;
   52147: out<=1;
   52148: out<=0;
   52149: out<=0;
   52150: out<=0;
   52151: out<=0;
   52152: out<=0;
   52153: out<=0;
   52154: out<=1;
   52155: out<=1;
   52156: out<=1;
   52157: out<=0;
   52158: out<=1;
   52159: out<=0;
   52160: out<=0;
   52161: out<=1;
   52162: out<=1;
   52163: out<=0;
   52164: out<=1;
   52165: out<=1;
   52166: out<=1;
   52167: out<=1;
   52168: out<=1;
   52169: out<=1;
   52170: out<=0;
   52171: out<=0;
   52172: out<=0;
   52173: out<=1;
   52174: out<=0;
   52175: out<=1;
   52176: out<=1;
   52177: out<=0;
   52178: out<=0;
   52179: out<=1;
   52180: out<=0;
   52181: out<=0;
   52182: out<=0;
   52183: out<=0;
   52184: out<=0;
   52185: out<=0;
   52186: out<=1;
   52187: out<=1;
   52188: out<=1;
   52189: out<=0;
   52190: out<=1;
   52191: out<=0;
   52192: out<=1;
   52193: out<=0;
   52194: out<=0;
   52195: out<=1;
   52196: out<=0;
   52197: out<=0;
   52198: out<=0;
   52199: out<=0;
   52200: out<=0;
   52201: out<=0;
   52202: out<=1;
   52203: out<=1;
   52204: out<=1;
   52205: out<=0;
   52206: out<=1;
   52207: out<=0;
   52208: out<=0;
   52209: out<=1;
   52210: out<=1;
   52211: out<=0;
   52212: out<=1;
   52213: out<=1;
   52214: out<=1;
   52215: out<=1;
   52216: out<=1;
   52217: out<=1;
   52218: out<=0;
   52219: out<=0;
   52220: out<=0;
   52221: out<=1;
   52222: out<=0;
   52223: out<=1;
   52224: out<=0;
   52225: out<=0;
   52226: out<=1;
   52227: out<=1;
   52228: out<=1;
   52229: out<=0;
   52230: out<=1;
   52231: out<=0;
   52232: out<=0;
   52233: out<=1;
   52234: out<=1;
   52235: out<=0;
   52236: out<=1;
   52237: out<=1;
   52238: out<=1;
   52239: out<=1;
   52240: out<=1;
   52241: out<=1;
   52242: out<=0;
   52243: out<=0;
   52244: out<=0;
   52245: out<=1;
   52246: out<=0;
   52247: out<=1;
   52248: out<=1;
   52249: out<=0;
   52250: out<=0;
   52251: out<=1;
   52252: out<=0;
   52253: out<=0;
   52254: out<=0;
   52255: out<=0;
   52256: out<=1;
   52257: out<=1;
   52258: out<=0;
   52259: out<=0;
   52260: out<=0;
   52261: out<=1;
   52262: out<=0;
   52263: out<=1;
   52264: out<=1;
   52265: out<=0;
   52266: out<=0;
   52267: out<=1;
   52268: out<=0;
   52269: out<=0;
   52270: out<=0;
   52271: out<=0;
   52272: out<=0;
   52273: out<=0;
   52274: out<=1;
   52275: out<=1;
   52276: out<=1;
   52277: out<=0;
   52278: out<=1;
   52279: out<=0;
   52280: out<=0;
   52281: out<=1;
   52282: out<=1;
   52283: out<=0;
   52284: out<=1;
   52285: out<=1;
   52286: out<=1;
   52287: out<=1;
   52288: out<=1;
   52289: out<=1;
   52290: out<=0;
   52291: out<=0;
   52292: out<=0;
   52293: out<=1;
   52294: out<=0;
   52295: out<=1;
   52296: out<=1;
   52297: out<=0;
   52298: out<=0;
   52299: out<=1;
   52300: out<=0;
   52301: out<=0;
   52302: out<=0;
   52303: out<=0;
   52304: out<=1;
   52305: out<=1;
   52306: out<=0;
   52307: out<=0;
   52308: out<=0;
   52309: out<=1;
   52310: out<=0;
   52311: out<=1;
   52312: out<=1;
   52313: out<=0;
   52314: out<=0;
   52315: out<=1;
   52316: out<=0;
   52317: out<=0;
   52318: out<=0;
   52319: out<=0;
   52320: out<=1;
   52321: out<=1;
   52322: out<=0;
   52323: out<=0;
   52324: out<=0;
   52325: out<=1;
   52326: out<=0;
   52327: out<=1;
   52328: out<=1;
   52329: out<=0;
   52330: out<=0;
   52331: out<=1;
   52332: out<=0;
   52333: out<=0;
   52334: out<=0;
   52335: out<=0;
   52336: out<=1;
   52337: out<=1;
   52338: out<=0;
   52339: out<=0;
   52340: out<=0;
   52341: out<=1;
   52342: out<=0;
   52343: out<=1;
   52344: out<=1;
   52345: out<=0;
   52346: out<=0;
   52347: out<=1;
   52348: out<=0;
   52349: out<=0;
   52350: out<=0;
   52351: out<=0;
   52352: out<=0;
   52353: out<=0;
   52354: out<=1;
   52355: out<=1;
   52356: out<=1;
   52357: out<=0;
   52358: out<=1;
   52359: out<=0;
   52360: out<=0;
   52361: out<=1;
   52362: out<=1;
   52363: out<=0;
   52364: out<=1;
   52365: out<=1;
   52366: out<=1;
   52367: out<=1;
   52368: out<=0;
   52369: out<=0;
   52370: out<=1;
   52371: out<=1;
   52372: out<=1;
   52373: out<=0;
   52374: out<=1;
   52375: out<=0;
   52376: out<=0;
   52377: out<=1;
   52378: out<=1;
   52379: out<=0;
   52380: out<=1;
   52381: out<=1;
   52382: out<=1;
   52383: out<=1;
   52384: out<=1;
   52385: out<=1;
   52386: out<=0;
   52387: out<=0;
   52388: out<=0;
   52389: out<=1;
   52390: out<=0;
   52391: out<=1;
   52392: out<=1;
   52393: out<=0;
   52394: out<=0;
   52395: out<=1;
   52396: out<=0;
   52397: out<=0;
   52398: out<=0;
   52399: out<=0;
   52400: out<=1;
   52401: out<=1;
   52402: out<=0;
   52403: out<=0;
   52404: out<=0;
   52405: out<=1;
   52406: out<=0;
   52407: out<=1;
   52408: out<=1;
   52409: out<=0;
   52410: out<=0;
   52411: out<=1;
   52412: out<=0;
   52413: out<=0;
   52414: out<=0;
   52415: out<=0;
   52416: out<=1;
   52417: out<=1;
   52418: out<=0;
   52419: out<=0;
   52420: out<=0;
   52421: out<=1;
   52422: out<=0;
   52423: out<=1;
   52424: out<=1;
   52425: out<=0;
   52426: out<=0;
   52427: out<=1;
   52428: out<=0;
   52429: out<=0;
   52430: out<=0;
   52431: out<=0;
   52432: out<=0;
   52433: out<=0;
   52434: out<=1;
   52435: out<=1;
   52436: out<=1;
   52437: out<=0;
   52438: out<=1;
   52439: out<=0;
   52440: out<=0;
   52441: out<=1;
   52442: out<=1;
   52443: out<=0;
   52444: out<=1;
   52445: out<=1;
   52446: out<=1;
   52447: out<=1;
   52448: out<=1;
   52449: out<=1;
   52450: out<=0;
   52451: out<=0;
   52452: out<=0;
   52453: out<=1;
   52454: out<=0;
   52455: out<=1;
   52456: out<=1;
   52457: out<=0;
   52458: out<=0;
   52459: out<=1;
   52460: out<=0;
   52461: out<=0;
   52462: out<=0;
   52463: out<=0;
   52464: out<=0;
   52465: out<=0;
   52466: out<=1;
   52467: out<=1;
   52468: out<=1;
   52469: out<=0;
   52470: out<=1;
   52471: out<=0;
   52472: out<=0;
   52473: out<=1;
   52474: out<=1;
   52475: out<=0;
   52476: out<=1;
   52477: out<=1;
   52478: out<=1;
   52479: out<=1;
   52480: out<=0;
   52481: out<=1;
   52482: out<=0;
   52483: out<=1;
   52484: out<=0;
   52485: out<=0;
   52486: out<=1;
   52487: out<=1;
   52488: out<=1;
   52489: out<=1;
   52490: out<=1;
   52491: out<=1;
   52492: out<=1;
   52493: out<=0;
   52494: out<=0;
   52495: out<=1;
   52496: out<=0;
   52497: out<=1;
   52498: out<=0;
   52499: out<=1;
   52500: out<=0;
   52501: out<=0;
   52502: out<=1;
   52503: out<=1;
   52504: out<=1;
   52505: out<=1;
   52506: out<=1;
   52507: out<=1;
   52508: out<=1;
   52509: out<=0;
   52510: out<=0;
   52511: out<=1;
   52512: out<=0;
   52513: out<=1;
   52514: out<=0;
   52515: out<=1;
   52516: out<=0;
   52517: out<=0;
   52518: out<=1;
   52519: out<=1;
   52520: out<=1;
   52521: out<=1;
   52522: out<=1;
   52523: out<=1;
   52524: out<=1;
   52525: out<=0;
   52526: out<=0;
   52527: out<=1;
   52528: out<=0;
   52529: out<=1;
   52530: out<=0;
   52531: out<=1;
   52532: out<=0;
   52533: out<=0;
   52534: out<=1;
   52535: out<=1;
   52536: out<=1;
   52537: out<=1;
   52538: out<=1;
   52539: out<=1;
   52540: out<=1;
   52541: out<=0;
   52542: out<=0;
   52543: out<=1;
   52544: out<=1;
   52545: out<=0;
   52546: out<=1;
   52547: out<=0;
   52548: out<=1;
   52549: out<=1;
   52550: out<=0;
   52551: out<=0;
   52552: out<=0;
   52553: out<=0;
   52554: out<=0;
   52555: out<=0;
   52556: out<=0;
   52557: out<=1;
   52558: out<=1;
   52559: out<=0;
   52560: out<=0;
   52561: out<=1;
   52562: out<=0;
   52563: out<=1;
   52564: out<=0;
   52565: out<=0;
   52566: out<=1;
   52567: out<=1;
   52568: out<=1;
   52569: out<=1;
   52570: out<=1;
   52571: out<=1;
   52572: out<=1;
   52573: out<=0;
   52574: out<=0;
   52575: out<=1;
   52576: out<=0;
   52577: out<=1;
   52578: out<=0;
   52579: out<=1;
   52580: out<=0;
   52581: out<=0;
   52582: out<=1;
   52583: out<=1;
   52584: out<=1;
   52585: out<=1;
   52586: out<=1;
   52587: out<=1;
   52588: out<=1;
   52589: out<=0;
   52590: out<=0;
   52591: out<=1;
   52592: out<=1;
   52593: out<=0;
   52594: out<=1;
   52595: out<=0;
   52596: out<=1;
   52597: out<=1;
   52598: out<=0;
   52599: out<=0;
   52600: out<=0;
   52601: out<=0;
   52602: out<=0;
   52603: out<=0;
   52604: out<=0;
   52605: out<=1;
   52606: out<=1;
   52607: out<=0;
   52608: out<=0;
   52609: out<=1;
   52610: out<=0;
   52611: out<=1;
   52612: out<=0;
   52613: out<=0;
   52614: out<=1;
   52615: out<=1;
   52616: out<=1;
   52617: out<=1;
   52618: out<=1;
   52619: out<=1;
   52620: out<=1;
   52621: out<=0;
   52622: out<=0;
   52623: out<=1;
   52624: out<=1;
   52625: out<=0;
   52626: out<=1;
   52627: out<=0;
   52628: out<=1;
   52629: out<=1;
   52630: out<=0;
   52631: out<=0;
   52632: out<=0;
   52633: out<=0;
   52634: out<=0;
   52635: out<=0;
   52636: out<=0;
   52637: out<=1;
   52638: out<=1;
   52639: out<=0;
   52640: out<=0;
   52641: out<=1;
   52642: out<=0;
   52643: out<=1;
   52644: out<=0;
   52645: out<=0;
   52646: out<=1;
   52647: out<=1;
   52648: out<=1;
   52649: out<=1;
   52650: out<=1;
   52651: out<=1;
   52652: out<=1;
   52653: out<=0;
   52654: out<=0;
   52655: out<=1;
   52656: out<=1;
   52657: out<=0;
   52658: out<=1;
   52659: out<=0;
   52660: out<=1;
   52661: out<=1;
   52662: out<=0;
   52663: out<=0;
   52664: out<=0;
   52665: out<=0;
   52666: out<=0;
   52667: out<=0;
   52668: out<=0;
   52669: out<=1;
   52670: out<=1;
   52671: out<=0;
   52672: out<=1;
   52673: out<=0;
   52674: out<=1;
   52675: out<=0;
   52676: out<=1;
   52677: out<=1;
   52678: out<=0;
   52679: out<=0;
   52680: out<=0;
   52681: out<=0;
   52682: out<=0;
   52683: out<=0;
   52684: out<=0;
   52685: out<=1;
   52686: out<=1;
   52687: out<=0;
   52688: out<=1;
   52689: out<=0;
   52690: out<=1;
   52691: out<=0;
   52692: out<=1;
   52693: out<=1;
   52694: out<=0;
   52695: out<=0;
   52696: out<=0;
   52697: out<=0;
   52698: out<=0;
   52699: out<=0;
   52700: out<=0;
   52701: out<=1;
   52702: out<=1;
   52703: out<=0;
   52704: out<=0;
   52705: out<=1;
   52706: out<=0;
   52707: out<=1;
   52708: out<=0;
   52709: out<=0;
   52710: out<=1;
   52711: out<=1;
   52712: out<=1;
   52713: out<=1;
   52714: out<=1;
   52715: out<=1;
   52716: out<=1;
   52717: out<=0;
   52718: out<=0;
   52719: out<=1;
   52720: out<=0;
   52721: out<=1;
   52722: out<=0;
   52723: out<=1;
   52724: out<=0;
   52725: out<=0;
   52726: out<=1;
   52727: out<=1;
   52728: out<=1;
   52729: out<=1;
   52730: out<=1;
   52731: out<=1;
   52732: out<=1;
   52733: out<=0;
   52734: out<=0;
   52735: out<=1;
   52736: out<=1;
   52737: out<=0;
   52738: out<=0;
   52739: out<=1;
   52740: out<=1;
   52741: out<=1;
   52742: out<=1;
   52743: out<=1;
   52744: out<=1;
   52745: out<=1;
   52746: out<=0;
   52747: out<=0;
   52748: out<=1;
   52749: out<=0;
   52750: out<=1;
   52751: out<=0;
   52752: out<=1;
   52753: out<=0;
   52754: out<=0;
   52755: out<=1;
   52756: out<=1;
   52757: out<=1;
   52758: out<=1;
   52759: out<=1;
   52760: out<=1;
   52761: out<=1;
   52762: out<=0;
   52763: out<=0;
   52764: out<=1;
   52765: out<=0;
   52766: out<=1;
   52767: out<=0;
   52768: out<=0;
   52769: out<=1;
   52770: out<=1;
   52771: out<=0;
   52772: out<=0;
   52773: out<=0;
   52774: out<=0;
   52775: out<=0;
   52776: out<=0;
   52777: out<=0;
   52778: out<=1;
   52779: out<=1;
   52780: out<=0;
   52781: out<=1;
   52782: out<=0;
   52783: out<=1;
   52784: out<=0;
   52785: out<=1;
   52786: out<=1;
   52787: out<=0;
   52788: out<=0;
   52789: out<=0;
   52790: out<=0;
   52791: out<=0;
   52792: out<=0;
   52793: out<=0;
   52794: out<=1;
   52795: out<=1;
   52796: out<=0;
   52797: out<=1;
   52798: out<=0;
   52799: out<=1;
   52800: out<=0;
   52801: out<=1;
   52802: out<=1;
   52803: out<=0;
   52804: out<=0;
   52805: out<=0;
   52806: out<=0;
   52807: out<=0;
   52808: out<=0;
   52809: out<=0;
   52810: out<=1;
   52811: out<=1;
   52812: out<=0;
   52813: out<=1;
   52814: out<=0;
   52815: out<=1;
   52816: out<=1;
   52817: out<=0;
   52818: out<=0;
   52819: out<=1;
   52820: out<=1;
   52821: out<=1;
   52822: out<=1;
   52823: out<=1;
   52824: out<=1;
   52825: out<=1;
   52826: out<=0;
   52827: out<=0;
   52828: out<=1;
   52829: out<=0;
   52830: out<=1;
   52831: out<=0;
   52832: out<=0;
   52833: out<=1;
   52834: out<=1;
   52835: out<=0;
   52836: out<=0;
   52837: out<=0;
   52838: out<=0;
   52839: out<=0;
   52840: out<=0;
   52841: out<=0;
   52842: out<=1;
   52843: out<=1;
   52844: out<=0;
   52845: out<=1;
   52846: out<=0;
   52847: out<=1;
   52848: out<=1;
   52849: out<=0;
   52850: out<=0;
   52851: out<=1;
   52852: out<=1;
   52853: out<=1;
   52854: out<=1;
   52855: out<=1;
   52856: out<=1;
   52857: out<=1;
   52858: out<=0;
   52859: out<=0;
   52860: out<=1;
   52861: out<=0;
   52862: out<=1;
   52863: out<=0;
   52864: out<=1;
   52865: out<=0;
   52866: out<=0;
   52867: out<=1;
   52868: out<=1;
   52869: out<=1;
   52870: out<=1;
   52871: out<=1;
   52872: out<=1;
   52873: out<=1;
   52874: out<=0;
   52875: out<=0;
   52876: out<=1;
   52877: out<=0;
   52878: out<=1;
   52879: out<=0;
   52880: out<=0;
   52881: out<=1;
   52882: out<=1;
   52883: out<=0;
   52884: out<=0;
   52885: out<=0;
   52886: out<=0;
   52887: out<=0;
   52888: out<=0;
   52889: out<=0;
   52890: out<=1;
   52891: out<=1;
   52892: out<=0;
   52893: out<=1;
   52894: out<=0;
   52895: out<=1;
   52896: out<=0;
   52897: out<=1;
   52898: out<=1;
   52899: out<=0;
   52900: out<=0;
   52901: out<=0;
   52902: out<=0;
   52903: out<=0;
   52904: out<=0;
   52905: out<=0;
   52906: out<=1;
   52907: out<=1;
   52908: out<=0;
   52909: out<=1;
   52910: out<=0;
   52911: out<=1;
   52912: out<=1;
   52913: out<=0;
   52914: out<=0;
   52915: out<=1;
   52916: out<=1;
   52917: out<=1;
   52918: out<=1;
   52919: out<=1;
   52920: out<=1;
   52921: out<=1;
   52922: out<=0;
   52923: out<=0;
   52924: out<=1;
   52925: out<=0;
   52926: out<=1;
   52927: out<=0;
   52928: out<=0;
   52929: out<=1;
   52930: out<=1;
   52931: out<=0;
   52932: out<=0;
   52933: out<=0;
   52934: out<=0;
   52935: out<=0;
   52936: out<=0;
   52937: out<=0;
   52938: out<=1;
   52939: out<=1;
   52940: out<=0;
   52941: out<=1;
   52942: out<=0;
   52943: out<=1;
   52944: out<=0;
   52945: out<=1;
   52946: out<=1;
   52947: out<=0;
   52948: out<=0;
   52949: out<=0;
   52950: out<=0;
   52951: out<=0;
   52952: out<=0;
   52953: out<=0;
   52954: out<=1;
   52955: out<=1;
   52956: out<=0;
   52957: out<=1;
   52958: out<=0;
   52959: out<=1;
   52960: out<=0;
   52961: out<=1;
   52962: out<=1;
   52963: out<=0;
   52964: out<=0;
   52965: out<=0;
   52966: out<=0;
   52967: out<=0;
   52968: out<=0;
   52969: out<=0;
   52970: out<=1;
   52971: out<=1;
   52972: out<=0;
   52973: out<=1;
   52974: out<=0;
   52975: out<=1;
   52976: out<=0;
   52977: out<=1;
   52978: out<=1;
   52979: out<=0;
   52980: out<=0;
   52981: out<=0;
   52982: out<=0;
   52983: out<=0;
   52984: out<=0;
   52985: out<=0;
   52986: out<=1;
   52987: out<=1;
   52988: out<=0;
   52989: out<=1;
   52990: out<=0;
   52991: out<=1;
   52992: out<=1;
   52993: out<=1;
   52994: out<=1;
   52995: out<=1;
   52996: out<=0;
   52997: out<=1;
   52998: out<=1;
   52999: out<=0;
   53000: out<=0;
   53001: out<=1;
   53002: out<=0;
   53003: out<=1;
   53004: out<=1;
   53005: out<=1;
   53006: out<=0;
   53007: out<=0;
   53008: out<=0;
   53009: out<=0;
   53010: out<=0;
   53011: out<=0;
   53012: out<=1;
   53013: out<=0;
   53014: out<=0;
   53015: out<=1;
   53016: out<=1;
   53017: out<=0;
   53018: out<=1;
   53019: out<=0;
   53020: out<=0;
   53021: out<=0;
   53022: out<=1;
   53023: out<=1;
   53024: out<=1;
   53025: out<=1;
   53026: out<=1;
   53027: out<=1;
   53028: out<=0;
   53029: out<=1;
   53030: out<=1;
   53031: out<=0;
   53032: out<=0;
   53033: out<=1;
   53034: out<=0;
   53035: out<=1;
   53036: out<=1;
   53037: out<=1;
   53038: out<=0;
   53039: out<=0;
   53040: out<=0;
   53041: out<=0;
   53042: out<=0;
   53043: out<=0;
   53044: out<=1;
   53045: out<=0;
   53046: out<=0;
   53047: out<=1;
   53048: out<=1;
   53049: out<=0;
   53050: out<=1;
   53051: out<=0;
   53052: out<=0;
   53053: out<=0;
   53054: out<=1;
   53055: out<=1;
   53056: out<=0;
   53057: out<=0;
   53058: out<=0;
   53059: out<=0;
   53060: out<=1;
   53061: out<=0;
   53062: out<=0;
   53063: out<=1;
   53064: out<=1;
   53065: out<=0;
   53066: out<=1;
   53067: out<=0;
   53068: out<=0;
   53069: out<=0;
   53070: out<=1;
   53071: out<=1;
   53072: out<=0;
   53073: out<=0;
   53074: out<=0;
   53075: out<=0;
   53076: out<=1;
   53077: out<=0;
   53078: out<=0;
   53079: out<=1;
   53080: out<=1;
   53081: out<=0;
   53082: out<=1;
   53083: out<=0;
   53084: out<=0;
   53085: out<=0;
   53086: out<=1;
   53087: out<=1;
   53088: out<=1;
   53089: out<=1;
   53090: out<=1;
   53091: out<=1;
   53092: out<=0;
   53093: out<=1;
   53094: out<=1;
   53095: out<=0;
   53096: out<=0;
   53097: out<=1;
   53098: out<=0;
   53099: out<=1;
   53100: out<=1;
   53101: out<=1;
   53102: out<=0;
   53103: out<=0;
   53104: out<=1;
   53105: out<=1;
   53106: out<=1;
   53107: out<=1;
   53108: out<=0;
   53109: out<=1;
   53110: out<=1;
   53111: out<=0;
   53112: out<=0;
   53113: out<=1;
   53114: out<=0;
   53115: out<=1;
   53116: out<=1;
   53117: out<=1;
   53118: out<=0;
   53119: out<=0;
   53120: out<=1;
   53121: out<=1;
   53122: out<=1;
   53123: out<=1;
   53124: out<=0;
   53125: out<=1;
   53126: out<=1;
   53127: out<=0;
   53128: out<=0;
   53129: out<=1;
   53130: out<=0;
   53131: out<=1;
   53132: out<=1;
   53133: out<=1;
   53134: out<=0;
   53135: out<=0;
   53136: out<=1;
   53137: out<=1;
   53138: out<=1;
   53139: out<=1;
   53140: out<=0;
   53141: out<=1;
   53142: out<=1;
   53143: out<=0;
   53144: out<=0;
   53145: out<=1;
   53146: out<=0;
   53147: out<=1;
   53148: out<=1;
   53149: out<=1;
   53150: out<=0;
   53151: out<=0;
   53152: out<=1;
   53153: out<=1;
   53154: out<=1;
   53155: out<=1;
   53156: out<=0;
   53157: out<=1;
   53158: out<=1;
   53159: out<=0;
   53160: out<=0;
   53161: out<=1;
   53162: out<=0;
   53163: out<=1;
   53164: out<=1;
   53165: out<=1;
   53166: out<=0;
   53167: out<=0;
   53168: out<=1;
   53169: out<=1;
   53170: out<=1;
   53171: out<=1;
   53172: out<=0;
   53173: out<=1;
   53174: out<=1;
   53175: out<=0;
   53176: out<=0;
   53177: out<=1;
   53178: out<=0;
   53179: out<=1;
   53180: out<=1;
   53181: out<=1;
   53182: out<=0;
   53183: out<=0;
   53184: out<=0;
   53185: out<=0;
   53186: out<=0;
   53187: out<=0;
   53188: out<=1;
   53189: out<=0;
   53190: out<=0;
   53191: out<=1;
   53192: out<=1;
   53193: out<=0;
   53194: out<=1;
   53195: out<=0;
   53196: out<=0;
   53197: out<=0;
   53198: out<=1;
   53199: out<=1;
   53200: out<=1;
   53201: out<=1;
   53202: out<=1;
   53203: out<=1;
   53204: out<=0;
   53205: out<=1;
   53206: out<=1;
   53207: out<=0;
   53208: out<=0;
   53209: out<=1;
   53210: out<=0;
   53211: out<=1;
   53212: out<=1;
   53213: out<=1;
   53214: out<=0;
   53215: out<=0;
   53216: out<=1;
   53217: out<=1;
   53218: out<=1;
   53219: out<=1;
   53220: out<=0;
   53221: out<=1;
   53222: out<=1;
   53223: out<=0;
   53224: out<=0;
   53225: out<=1;
   53226: out<=0;
   53227: out<=1;
   53228: out<=1;
   53229: out<=1;
   53230: out<=0;
   53231: out<=0;
   53232: out<=0;
   53233: out<=0;
   53234: out<=0;
   53235: out<=0;
   53236: out<=1;
   53237: out<=0;
   53238: out<=0;
   53239: out<=1;
   53240: out<=1;
   53241: out<=0;
   53242: out<=1;
   53243: out<=0;
   53244: out<=0;
   53245: out<=0;
   53246: out<=1;
   53247: out<=1;
   53248: out<=0;
   53249: out<=1;
   53250: out<=1;
   53251: out<=0;
   53252: out<=1;
   53253: out<=1;
   53254: out<=1;
   53255: out<=1;
   53256: out<=0;
   53257: out<=0;
   53258: out<=1;
   53259: out<=1;
   53260: out<=1;
   53261: out<=0;
   53262: out<=1;
   53263: out<=0;
   53264: out<=0;
   53265: out<=1;
   53266: out<=1;
   53267: out<=0;
   53268: out<=1;
   53269: out<=1;
   53270: out<=1;
   53271: out<=1;
   53272: out<=0;
   53273: out<=0;
   53274: out<=1;
   53275: out<=1;
   53276: out<=1;
   53277: out<=0;
   53278: out<=1;
   53279: out<=0;
   53280: out<=0;
   53281: out<=1;
   53282: out<=1;
   53283: out<=0;
   53284: out<=1;
   53285: out<=1;
   53286: out<=1;
   53287: out<=1;
   53288: out<=0;
   53289: out<=0;
   53290: out<=1;
   53291: out<=1;
   53292: out<=1;
   53293: out<=0;
   53294: out<=1;
   53295: out<=0;
   53296: out<=0;
   53297: out<=1;
   53298: out<=1;
   53299: out<=0;
   53300: out<=1;
   53301: out<=1;
   53302: out<=1;
   53303: out<=1;
   53304: out<=0;
   53305: out<=0;
   53306: out<=1;
   53307: out<=1;
   53308: out<=1;
   53309: out<=0;
   53310: out<=1;
   53311: out<=0;
   53312: out<=0;
   53313: out<=1;
   53314: out<=1;
   53315: out<=0;
   53316: out<=1;
   53317: out<=1;
   53318: out<=1;
   53319: out<=1;
   53320: out<=0;
   53321: out<=0;
   53322: out<=1;
   53323: out<=1;
   53324: out<=1;
   53325: out<=0;
   53326: out<=1;
   53327: out<=0;
   53328: out<=1;
   53329: out<=0;
   53330: out<=0;
   53331: out<=1;
   53332: out<=0;
   53333: out<=0;
   53334: out<=0;
   53335: out<=0;
   53336: out<=1;
   53337: out<=1;
   53338: out<=0;
   53339: out<=0;
   53340: out<=0;
   53341: out<=1;
   53342: out<=0;
   53343: out<=1;
   53344: out<=1;
   53345: out<=0;
   53346: out<=0;
   53347: out<=1;
   53348: out<=0;
   53349: out<=0;
   53350: out<=0;
   53351: out<=0;
   53352: out<=1;
   53353: out<=1;
   53354: out<=0;
   53355: out<=0;
   53356: out<=0;
   53357: out<=1;
   53358: out<=0;
   53359: out<=1;
   53360: out<=0;
   53361: out<=1;
   53362: out<=1;
   53363: out<=0;
   53364: out<=1;
   53365: out<=1;
   53366: out<=1;
   53367: out<=1;
   53368: out<=0;
   53369: out<=0;
   53370: out<=1;
   53371: out<=1;
   53372: out<=1;
   53373: out<=0;
   53374: out<=1;
   53375: out<=0;
   53376: out<=1;
   53377: out<=0;
   53378: out<=0;
   53379: out<=1;
   53380: out<=0;
   53381: out<=0;
   53382: out<=0;
   53383: out<=0;
   53384: out<=1;
   53385: out<=1;
   53386: out<=0;
   53387: out<=0;
   53388: out<=0;
   53389: out<=1;
   53390: out<=0;
   53391: out<=1;
   53392: out<=0;
   53393: out<=1;
   53394: out<=1;
   53395: out<=0;
   53396: out<=1;
   53397: out<=1;
   53398: out<=1;
   53399: out<=1;
   53400: out<=0;
   53401: out<=0;
   53402: out<=1;
   53403: out<=1;
   53404: out<=1;
   53405: out<=0;
   53406: out<=1;
   53407: out<=0;
   53408: out<=1;
   53409: out<=0;
   53410: out<=0;
   53411: out<=1;
   53412: out<=0;
   53413: out<=0;
   53414: out<=0;
   53415: out<=0;
   53416: out<=1;
   53417: out<=1;
   53418: out<=0;
   53419: out<=0;
   53420: out<=0;
   53421: out<=1;
   53422: out<=0;
   53423: out<=1;
   53424: out<=0;
   53425: out<=1;
   53426: out<=1;
   53427: out<=0;
   53428: out<=1;
   53429: out<=1;
   53430: out<=1;
   53431: out<=1;
   53432: out<=0;
   53433: out<=0;
   53434: out<=1;
   53435: out<=1;
   53436: out<=1;
   53437: out<=0;
   53438: out<=1;
   53439: out<=0;
   53440: out<=1;
   53441: out<=0;
   53442: out<=0;
   53443: out<=1;
   53444: out<=0;
   53445: out<=0;
   53446: out<=0;
   53447: out<=0;
   53448: out<=1;
   53449: out<=1;
   53450: out<=0;
   53451: out<=0;
   53452: out<=0;
   53453: out<=1;
   53454: out<=0;
   53455: out<=1;
   53456: out<=1;
   53457: out<=0;
   53458: out<=0;
   53459: out<=1;
   53460: out<=0;
   53461: out<=0;
   53462: out<=0;
   53463: out<=0;
   53464: out<=1;
   53465: out<=1;
   53466: out<=0;
   53467: out<=0;
   53468: out<=0;
   53469: out<=1;
   53470: out<=0;
   53471: out<=1;
   53472: out<=0;
   53473: out<=1;
   53474: out<=1;
   53475: out<=0;
   53476: out<=1;
   53477: out<=1;
   53478: out<=1;
   53479: out<=1;
   53480: out<=0;
   53481: out<=0;
   53482: out<=1;
   53483: out<=1;
   53484: out<=1;
   53485: out<=0;
   53486: out<=1;
   53487: out<=0;
   53488: out<=0;
   53489: out<=1;
   53490: out<=1;
   53491: out<=0;
   53492: out<=1;
   53493: out<=1;
   53494: out<=1;
   53495: out<=1;
   53496: out<=0;
   53497: out<=0;
   53498: out<=1;
   53499: out<=1;
   53500: out<=1;
   53501: out<=0;
   53502: out<=1;
   53503: out<=0;
   53504: out<=0;
   53505: out<=0;
   53506: out<=0;
   53507: out<=0;
   53508: out<=0;
   53509: out<=1;
   53510: out<=1;
   53511: out<=0;
   53512: out<=1;
   53513: out<=0;
   53514: out<=1;
   53515: out<=0;
   53516: out<=1;
   53517: out<=1;
   53518: out<=0;
   53519: out<=0;
   53520: out<=1;
   53521: out<=1;
   53522: out<=1;
   53523: out<=1;
   53524: out<=1;
   53525: out<=0;
   53526: out<=0;
   53527: out<=1;
   53528: out<=0;
   53529: out<=1;
   53530: out<=0;
   53531: out<=1;
   53532: out<=0;
   53533: out<=0;
   53534: out<=1;
   53535: out<=1;
   53536: out<=1;
   53537: out<=1;
   53538: out<=1;
   53539: out<=1;
   53540: out<=1;
   53541: out<=0;
   53542: out<=0;
   53543: out<=1;
   53544: out<=0;
   53545: out<=1;
   53546: out<=0;
   53547: out<=1;
   53548: out<=0;
   53549: out<=0;
   53550: out<=1;
   53551: out<=1;
   53552: out<=0;
   53553: out<=0;
   53554: out<=0;
   53555: out<=0;
   53556: out<=0;
   53557: out<=1;
   53558: out<=1;
   53559: out<=0;
   53560: out<=1;
   53561: out<=0;
   53562: out<=1;
   53563: out<=0;
   53564: out<=1;
   53565: out<=1;
   53566: out<=0;
   53567: out<=0;
   53568: out<=0;
   53569: out<=0;
   53570: out<=0;
   53571: out<=0;
   53572: out<=0;
   53573: out<=1;
   53574: out<=1;
   53575: out<=0;
   53576: out<=1;
   53577: out<=0;
   53578: out<=1;
   53579: out<=0;
   53580: out<=1;
   53581: out<=1;
   53582: out<=0;
   53583: out<=0;
   53584: out<=0;
   53585: out<=0;
   53586: out<=0;
   53587: out<=0;
   53588: out<=0;
   53589: out<=1;
   53590: out<=1;
   53591: out<=0;
   53592: out<=1;
   53593: out<=0;
   53594: out<=1;
   53595: out<=0;
   53596: out<=1;
   53597: out<=1;
   53598: out<=0;
   53599: out<=0;
   53600: out<=0;
   53601: out<=0;
   53602: out<=0;
   53603: out<=0;
   53604: out<=0;
   53605: out<=1;
   53606: out<=1;
   53607: out<=0;
   53608: out<=1;
   53609: out<=0;
   53610: out<=1;
   53611: out<=0;
   53612: out<=1;
   53613: out<=1;
   53614: out<=0;
   53615: out<=0;
   53616: out<=0;
   53617: out<=0;
   53618: out<=0;
   53619: out<=0;
   53620: out<=0;
   53621: out<=1;
   53622: out<=1;
   53623: out<=0;
   53624: out<=1;
   53625: out<=0;
   53626: out<=1;
   53627: out<=0;
   53628: out<=1;
   53629: out<=1;
   53630: out<=0;
   53631: out<=0;
   53632: out<=1;
   53633: out<=1;
   53634: out<=1;
   53635: out<=1;
   53636: out<=1;
   53637: out<=0;
   53638: out<=0;
   53639: out<=1;
   53640: out<=0;
   53641: out<=1;
   53642: out<=0;
   53643: out<=1;
   53644: out<=0;
   53645: out<=0;
   53646: out<=1;
   53647: out<=1;
   53648: out<=1;
   53649: out<=1;
   53650: out<=1;
   53651: out<=1;
   53652: out<=1;
   53653: out<=0;
   53654: out<=0;
   53655: out<=1;
   53656: out<=0;
   53657: out<=1;
   53658: out<=0;
   53659: out<=1;
   53660: out<=0;
   53661: out<=0;
   53662: out<=1;
   53663: out<=1;
   53664: out<=0;
   53665: out<=0;
   53666: out<=0;
   53667: out<=0;
   53668: out<=0;
   53669: out<=1;
   53670: out<=1;
   53671: out<=0;
   53672: out<=1;
   53673: out<=0;
   53674: out<=1;
   53675: out<=0;
   53676: out<=1;
   53677: out<=1;
   53678: out<=0;
   53679: out<=0;
   53680: out<=0;
   53681: out<=0;
   53682: out<=0;
   53683: out<=0;
   53684: out<=0;
   53685: out<=1;
   53686: out<=1;
   53687: out<=0;
   53688: out<=1;
   53689: out<=0;
   53690: out<=1;
   53691: out<=0;
   53692: out<=1;
   53693: out<=1;
   53694: out<=0;
   53695: out<=0;
   53696: out<=1;
   53697: out<=1;
   53698: out<=1;
   53699: out<=1;
   53700: out<=1;
   53701: out<=0;
   53702: out<=0;
   53703: out<=1;
   53704: out<=0;
   53705: out<=1;
   53706: out<=0;
   53707: out<=1;
   53708: out<=0;
   53709: out<=0;
   53710: out<=1;
   53711: out<=1;
   53712: out<=0;
   53713: out<=0;
   53714: out<=0;
   53715: out<=0;
   53716: out<=0;
   53717: out<=1;
   53718: out<=1;
   53719: out<=0;
   53720: out<=1;
   53721: out<=0;
   53722: out<=1;
   53723: out<=0;
   53724: out<=1;
   53725: out<=1;
   53726: out<=0;
   53727: out<=0;
   53728: out<=1;
   53729: out<=1;
   53730: out<=1;
   53731: out<=1;
   53732: out<=1;
   53733: out<=0;
   53734: out<=0;
   53735: out<=1;
   53736: out<=0;
   53737: out<=1;
   53738: out<=0;
   53739: out<=1;
   53740: out<=0;
   53741: out<=0;
   53742: out<=1;
   53743: out<=1;
   53744: out<=0;
   53745: out<=0;
   53746: out<=0;
   53747: out<=0;
   53748: out<=0;
   53749: out<=1;
   53750: out<=1;
   53751: out<=0;
   53752: out<=1;
   53753: out<=0;
   53754: out<=1;
   53755: out<=0;
   53756: out<=1;
   53757: out<=1;
   53758: out<=0;
   53759: out<=0;
   53760: out<=0;
   53761: out<=0;
   53762: out<=1;
   53763: out<=1;
   53764: out<=0;
   53765: out<=1;
   53766: out<=0;
   53767: out<=1;
   53768: out<=0;
   53769: out<=1;
   53770: out<=1;
   53771: out<=0;
   53772: out<=0;
   53773: out<=0;
   53774: out<=0;
   53775: out<=0;
   53776: out<=1;
   53777: out<=1;
   53778: out<=0;
   53779: out<=0;
   53780: out<=1;
   53781: out<=0;
   53782: out<=1;
   53783: out<=0;
   53784: out<=1;
   53785: out<=0;
   53786: out<=0;
   53787: out<=1;
   53788: out<=1;
   53789: out<=1;
   53790: out<=1;
   53791: out<=1;
   53792: out<=0;
   53793: out<=0;
   53794: out<=1;
   53795: out<=1;
   53796: out<=0;
   53797: out<=1;
   53798: out<=0;
   53799: out<=1;
   53800: out<=0;
   53801: out<=1;
   53802: out<=1;
   53803: out<=0;
   53804: out<=0;
   53805: out<=0;
   53806: out<=0;
   53807: out<=0;
   53808: out<=1;
   53809: out<=1;
   53810: out<=0;
   53811: out<=0;
   53812: out<=1;
   53813: out<=0;
   53814: out<=1;
   53815: out<=0;
   53816: out<=1;
   53817: out<=0;
   53818: out<=0;
   53819: out<=1;
   53820: out<=1;
   53821: out<=1;
   53822: out<=1;
   53823: out<=1;
   53824: out<=0;
   53825: out<=0;
   53826: out<=1;
   53827: out<=1;
   53828: out<=0;
   53829: out<=1;
   53830: out<=0;
   53831: out<=1;
   53832: out<=0;
   53833: out<=1;
   53834: out<=1;
   53835: out<=0;
   53836: out<=0;
   53837: out<=0;
   53838: out<=0;
   53839: out<=0;
   53840: out<=0;
   53841: out<=0;
   53842: out<=1;
   53843: out<=1;
   53844: out<=0;
   53845: out<=1;
   53846: out<=0;
   53847: out<=1;
   53848: out<=0;
   53849: out<=1;
   53850: out<=1;
   53851: out<=0;
   53852: out<=0;
   53853: out<=0;
   53854: out<=0;
   53855: out<=0;
   53856: out<=1;
   53857: out<=1;
   53858: out<=0;
   53859: out<=0;
   53860: out<=1;
   53861: out<=0;
   53862: out<=1;
   53863: out<=0;
   53864: out<=1;
   53865: out<=0;
   53866: out<=0;
   53867: out<=1;
   53868: out<=1;
   53869: out<=1;
   53870: out<=1;
   53871: out<=1;
   53872: out<=1;
   53873: out<=1;
   53874: out<=0;
   53875: out<=0;
   53876: out<=1;
   53877: out<=0;
   53878: out<=1;
   53879: out<=0;
   53880: out<=1;
   53881: out<=0;
   53882: out<=0;
   53883: out<=1;
   53884: out<=1;
   53885: out<=1;
   53886: out<=1;
   53887: out<=1;
   53888: out<=1;
   53889: out<=1;
   53890: out<=0;
   53891: out<=0;
   53892: out<=1;
   53893: out<=0;
   53894: out<=1;
   53895: out<=0;
   53896: out<=1;
   53897: out<=0;
   53898: out<=0;
   53899: out<=1;
   53900: out<=1;
   53901: out<=1;
   53902: out<=1;
   53903: out<=1;
   53904: out<=1;
   53905: out<=1;
   53906: out<=0;
   53907: out<=0;
   53908: out<=1;
   53909: out<=0;
   53910: out<=1;
   53911: out<=0;
   53912: out<=1;
   53913: out<=0;
   53914: out<=0;
   53915: out<=1;
   53916: out<=1;
   53917: out<=1;
   53918: out<=1;
   53919: out<=1;
   53920: out<=1;
   53921: out<=1;
   53922: out<=0;
   53923: out<=0;
   53924: out<=1;
   53925: out<=0;
   53926: out<=1;
   53927: out<=0;
   53928: out<=1;
   53929: out<=0;
   53930: out<=0;
   53931: out<=1;
   53932: out<=1;
   53933: out<=1;
   53934: out<=1;
   53935: out<=1;
   53936: out<=1;
   53937: out<=1;
   53938: out<=0;
   53939: out<=0;
   53940: out<=1;
   53941: out<=0;
   53942: out<=1;
   53943: out<=0;
   53944: out<=1;
   53945: out<=0;
   53946: out<=0;
   53947: out<=1;
   53948: out<=1;
   53949: out<=1;
   53950: out<=1;
   53951: out<=1;
   53952: out<=1;
   53953: out<=1;
   53954: out<=0;
   53955: out<=0;
   53956: out<=1;
   53957: out<=0;
   53958: out<=1;
   53959: out<=0;
   53960: out<=1;
   53961: out<=0;
   53962: out<=0;
   53963: out<=1;
   53964: out<=1;
   53965: out<=1;
   53966: out<=1;
   53967: out<=1;
   53968: out<=0;
   53969: out<=0;
   53970: out<=1;
   53971: out<=1;
   53972: out<=0;
   53973: out<=1;
   53974: out<=0;
   53975: out<=1;
   53976: out<=0;
   53977: out<=1;
   53978: out<=1;
   53979: out<=0;
   53980: out<=0;
   53981: out<=0;
   53982: out<=0;
   53983: out<=0;
   53984: out<=0;
   53985: out<=0;
   53986: out<=1;
   53987: out<=1;
   53988: out<=0;
   53989: out<=1;
   53990: out<=0;
   53991: out<=1;
   53992: out<=0;
   53993: out<=1;
   53994: out<=1;
   53995: out<=0;
   53996: out<=0;
   53997: out<=0;
   53998: out<=0;
   53999: out<=0;
   54000: out<=1;
   54001: out<=1;
   54002: out<=0;
   54003: out<=0;
   54004: out<=1;
   54005: out<=0;
   54006: out<=1;
   54007: out<=0;
   54008: out<=1;
   54009: out<=0;
   54010: out<=0;
   54011: out<=1;
   54012: out<=1;
   54013: out<=1;
   54014: out<=1;
   54015: out<=1;
   54016: out<=0;
   54017: out<=1;
   54018: out<=0;
   54019: out<=1;
   54020: out<=1;
   54021: out<=1;
   54022: out<=0;
   54023: out<=0;
   54024: out<=1;
   54025: out<=1;
   54026: out<=1;
   54027: out<=1;
   54028: out<=0;
   54029: out<=1;
   54030: out<=1;
   54031: out<=0;
   54032: out<=0;
   54033: out<=1;
   54034: out<=0;
   54035: out<=1;
   54036: out<=1;
   54037: out<=1;
   54038: out<=0;
   54039: out<=0;
   54040: out<=1;
   54041: out<=1;
   54042: out<=1;
   54043: out<=1;
   54044: out<=0;
   54045: out<=1;
   54046: out<=1;
   54047: out<=0;
   54048: out<=1;
   54049: out<=0;
   54050: out<=1;
   54051: out<=0;
   54052: out<=0;
   54053: out<=0;
   54054: out<=1;
   54055: out<=1;
   54056: out<=0;
   54057: out<=0;
   54058: out<=0;
   54059: out<=0;
   54060: out<=1;
   54061: out<=0;
   54062: out<=0;
   54063: out<=1;
   54064: out<=1;
   54065: out<=0;
   54066: out<=1;
   54067: out<=0;
   54068: out<=0;
   54069: out<=0;
   54070: out<=1;
   54071: out<=1;
   54072: out<=0;
   54073: out<=0;
   54074: out<=0;
   54075: out<=0;
   54076: out<=1;
   54077: out<=0;
   54078: out<=0;
   54079: out<=1;
   54080: out<=0;
   54081: out<=1;
   54082: out<=0;
   54083: out<=1;
   54084: out<=1;
   54085: out<=1;
   54086: out<=0;
   54087: out<=0;
   54088: out<=1;
   54089: out<=1;
   54090: out<=1;
   54091: out<=1;
   54092: out<=0;
   54093: out<=1;
   54094: out<=1;
   54095: out<=0;
   54096: out<=1;
   54097: out<=0;
   54098: out<=1;
   54099: out<=0;
   54100: out<=0;
   54101: out<=0;
   54102: out<=1;
   54103: out<=1;
   54104: out<=0;
   54105: out<=0;
   54106: out<=0;
   54107: out<=0;
   54108: out<=1;
   54109: out<=0;
   54110: out<=0;
   54111: out<=1;
   54112: out<=0;
   54113: out<=1;
   54114: out<=0;
   54115: out<=1;
   54116: out<=1;
   54117: out<=1;
   54118: out<=0;
   54119: out<=0;
   54120: out<=1;
   54121: out<=1;
   54122: out<=1;
   54123: out<=1;
   54124: out<=0;
   54125: out<=1;
   54126: out<=1;
   54127: out<=0;
   54128: out<=1;
   54129: out<=0;
   54130: out<=1;
   54131: out<=0;
   54132: out<=0;
   54133: out<=0;
   54134: out<=1;
   54135: out<=1;
   54136: out<=0;
   54137: out<=0;
   54138: out<=0;
   54139: out<=0;
   54140: out<=1;
   54141: out<=0;
   54142: out<=0;
   54143: out<=1;
   54144: out<=1;
   54145: out<=0;
   54146: out<=1;
   54147: out<=0;
   54148: out<=0;
   54149: out<=0;
   54150: out<=1;
   54151: out<=1;
   54152: out<=0;
   54153: out<=0;
   54154: out<=0;
   54155: out<=0;
   54156: out<=1;
   54157: out<=0;
   54158: out<=0;
   54159: out<=1;
   54160: out<=0;
   54161: out<=1;
   54162: out<=0;
   54163: out<=1;
   54164: out<=1;
   54165: out<=1;
   54166: out<=0;
   54167: out<=0;
   54168: out<=1;
   54169: out<=1;
   54170: out<=1;
   54171: out<=1;
   54172: out<=0;
   54173: out<=1;
   54174: out<=1;
   54175: out<=0;
   54176: out<=0;
   54177: out<=1;
   54178: out<=0;
   54179: out<=1;
   54180: out<=1;
   54181: out<=1;
   54182: out<=0;
   54183: out<=0;
   54184: out<=1;
   54185: out<=1;
   54186: out<=1;
   54187: out<=1;
   54188: out<=0;
   54189: out<=1;
   54190: out<=1;
   54191: out<=0;
   54192: out<=1;
   54193: out<=0;
   54194: out<=1;
   54195: out<=0;
   54196: out<=0;
   54197: out<=0;
   54198: out<=1;
   54199: out<=1;
   54200: out<=0;
   54201: out<=0;
   54202: out<=0;
   54203: out<=0;
   54204: out<=1;
   54205: out<=0;
   54206: out<=0;
   54207: out<=1;
   54208: out<=1;
   54209: out<=0;
   54210: out<=1;
   54211: out<=0;
   54212: out<=0;
   54213: out<=0;
   54214: out<=1;
   54215: out<=1;
   54216: out<=0;
   54217: out<=0;
   54218: out<=0;
   54219: out<=0;
   54220: out<=1;
   54221: out<=0;
   54222: out<=0;
   54223: out<=1;
   54224: out<=1;
   54225: out<=0;
   54226: out<=1;
   54227: out<=0;
   54228: out<=0;
   54229: out<=0;
   54230: out<=1;
   54231: out<=1;
   54232: out<=0;
   54233: out<=0;
   54234: out<=0;
   54235: out<=0;
   54236: out<=1;
   54237: out<=0;
   54238: out<=0;
   54239: out<=1;
   54240: out<=1;
   54241: out<=0;
   54242: out<=1;
   54243: out<=0;
   54244: out<=0;
   54245: out<=0;
   54246: out<=1;
   54247: out<=1;
   54248: out<=0;
   54249: out<=0;
   54250: out<=0;
   54251: out<=0;
   54252: out<=1;
   54253: out<=0;
   54254: out<=0;
   54255: out<=1;
   54256: out<=1;
   54257: out<=0;
   54258: out<=1;
   54259: out<=0;
   54260: out<=0;
   54261: out<=0;
   54262: out<=1;
   54263: out<=1;
   54264: out<=0;
   54265: out<=0;
   54266: out<=0;
   54267: out<=0;
   54268: out<=1;
   54269: out<=0;
   54270: out<=0;
   54271: out<=1;
   54272: out<=0;
   54273: out<=0;
   54274: out<=0;
   54275: out<=0;
   54276: out<=1;
   54277: out<=0;
   54278: out<=0;
   54279: out<=1;
   54280: out<=0;
   54281: out<=1;
   54282: out<=0;
   54283: out<=1;
   54284: out<=1;
   54285: out<=1;
   54286: out<=0;
   54287: out<=0;
   54288: out<=0;
   54289: out<=0;
   54290: out<=0;
   54291: out<=0;
   54292: out<=1;
   54293: out<=0;
   54294: out<=0;
   54295: out<=1;
   54296: out<=0;
   54297: out<=1;
   54298: out<=0;
   54299: out<=1;
   54300: out<=1;
   54301: out<=1;
   54302: out<=0;
   54303: out<=0;
   54304: out<=0;
   54305: out<=0;
   54306: out<=0;
   54307: out<=0;
   54308: out<=1;
   54309: out<=0;
   54310: out<=0;
   54311: out<=1;
   54312: out<=0;
   54313: out<=1;
   54314: out<=0;
   54315: out<=1;
   54316: out<=1;
   54317: out<=1;
   54318: out<=0;
   54319: out<=0;
   54320: out<=0;
   54321: out<=0;
   54322: out<=0;
   54323: out<=0;
   54324: out<=1;
   54325: out<=0;
   54326: out<=0;
   54327: out<=1;
   54328: out<=0;
   54329: out<=1;
   54330: out<=0;
   54331: out<=1;
   54332: out<=1;
   54333: out<=1;
   54334: out<=0;
   54335: out<=0;
   54336: out<=0;
   54337: out<=0;
   54338: out<=0;
   54339: out<=0;
   54340: out<=1;
   54341: out<=0;
   54342: out<=0;
   54343: out<=1;
   54344: out<=0;
   54345: out<=1;
   54346: out<=0;
   54347: out<=1;
   54348: out<=1;
   54349: out<=1;
   54350: out<=0;
   54351: out<=0;
   54352: out<=1;
   54353: out<=1;
   54354: out<=1;
   54355: out<=1;
   54356: out<=0;
   54357: out<=1;
   54358: out<=1;
   54359: out<=0;
   54360: out<=1;
   54361: out<=0;
   54362: out<=1;
   54363: out<=0;
   54364: out<=0;
   54365: out<=0;
   54366: out<=1;
   54367: out<=1;
   54368: out<=1;
   54369: out<=1;
   54370: out<=1;
   54371: out<=1;
   54372: out<=0;
   54373: out<=1;
   54374: out<=1;
   54375: out<=0;
   54376: out<=1;
   54377: out<=0;
   54378: out<=1;
   54379: out<=0;
   54380: out<=0;
   54381: out<=0;
   54382: out<=1;
   54383: out<=1;
   54384: out<=0;
   54385: out<=0;
   54386: out<=0;
   54387: out<=0;
   54388: out<=1;
   54389: out<=0;
   54390: out<=0;
   54391: out<=1;
   54392: out<=0;
   54393: out<=1;
   54394: out<=0;
   54395: out<=1;
   54396: out<=1;
   54397: out<=1;
   54398: out<=0;
   54399: out<=0;
   54400: out<=1;
   54401: out<=1;
   54402: out<=1;
   54403: out<=1;
   54404: out<=0;
   54405: out<=1;
   54406: out<=1;
   54407: out<=0;
   54408: out<=1;
   54409: out<=0;
   54410: out<=1;
   54411: out<=0;
   54412: out<=0;
   54413: out<=0;
   54414: out<=1;
   54415: out<=1;
   54416: out<=0;
   54417: out<=0;
   54418: out<=0;
   54419: out<=0;
   54420: out<=1;
   54421: out<=0;
   54422: out<=0;
   54423: out<=1;
   54424: out<=0;
   54425: out<=1;
   54426: out<=0;
   54427: out<=1;
   54428: out<=1;
   54429: out<=1;
   54430: out<=0;
   54431: out<=0;
   54432: out<=1;
   54433: out<=1;
   54434: out<=1;
   54435: out<=1;
   54436: out<=0;
   54437: out<=1;
   54438: out<=1;
   54439: out<=0;
   54440: out<=1;
   54441: out<=0;
   54442: out<=1;
   54443: out<=0;
   54444: out<=0;
   54445: out<=0;
   54446: out<=1;
   54447: out<=1;
   54448: out<=0;
   54449: out<=0;
   54450: out<=0;
   54451: out<=0;
   54452: out<=1;
   54453: out<=0;
   54454: out<=0;
   54455: out<=1;
   54456: out<=0;
   54457: out<=1;
   54458: out<=0;
   54459: out<=1;
   54460: out<=1;
   54461: out<=1;
   54462: out<=0;
   54463: out<=0;
   54464: out<=1;
   54465: out<=1;
   54466: out<=1;
   54467: out<=1;
   54468: out<=0;
   54469: out<=1;
   54470: out<=1;
   54471: out<=0;
   54472: out<=1;
   54473: out<=0;
   54474: out<=1;
   54475: out<=0;
   54476: out<=0;
   54477: out<=0;
   54478: out<=1;
   54479: out<=1;
   54480: out<=1;
   54481: out<=1;
   54482: out<=1;
   54483: out<=1;
   54484: out<=0;
   54485: out<=1;
   54486: out<=1;
   54487: out<=0;
   54488: out<=1;
   54489: out<=0;
   54490: out<=1;
   54491: out<=0;
   54492: out<=0;
   54493: out<=0;
   54494: out<=1;
   54495: out<=1;
   54496: out<=0;
   54497: out<=0;
   54498: out<=0;
   54499: out<=0;
   54500: out<=1;
   54501: out<=0;
   54502: out<=0;
   54503: out<=1;
   54504: out<=0;
   54505: out<=1;
   54506: out<=0;
   54507: out<=1;
   54508: out<=1;
   54509: out<=1;
   54510: out<=0;
   54511: out<=0;
   54512: out<=0;
   54513: out<=0;
   54514: out<=0;
   54515: out<=0;
   54516: out<=1;
   54517: out<=0;
   54518: out<=0;
   54519: out<=1;
   54520: out<=0;
   54521: out<=1;
   54522: out<=0;
   54523: out<=1;
   54524: out<=1;
   54525: out<=1;
   54526: out<=0;
   54527: out<=0;
   54528: out<=1;
   54529: out<=0;
   54530: out<=0;
   54531: out<=1;
   54532: out<=1;
   54533: out<=1;
   54534: out<=1;
   54535: out<=1;
   54536: out<=0;
   54537: out<=0;
   54538: out<=1;
   54539: out<=1;
   54540: out<=0;
   54541: out<=1;
   54542: out<=0;
   54543: out<=1;
   54544: out<=0;
   54545: out<=1;
   54546: out<=1;
   54547: out<=0;
   54548: out<=0;
   54549: out<=0;
   54550: out<=0;
   54551: out<=0;
   54552: out<=1;
   54553: out<=1;
   54554: out<=0;
   54555: out<=0;
   54556: out<=1;
   54557: out<=0;
   54558: out<=1;
   54559: out<=0;
   54560: out<=0;
   54561: out<=1;
   54562: out<=1;
   54563: out<=0;
   54564: out<=0;
   54565: out<=0;
   54566: out<=0;
   54567: out<=0;
   54568: out<=1;
   54569: out<=1;
   54570: out<=0;
   54571: out<=0;
   54572: out<=1;
   54573: out<=0;
   54574: out<=1;
   54575: out<=0;
   54576: out<=1;
   54577: out<=0;
   54578: out<=0;
   54579: out<=1;
   54580: out<=1;
   54581: out<=1;
   54582: out<=1;
   54583: out<=1;
   54584: out<=0;
   54585: out<=0;
   54586: out<=1;
   54587: out<=1;
   54588: out<=0;
   54589: out<=1;
   54590: out<=0;
   54591: out<=1;
   54592: out<=1;
   54593: out<=0;
   54594: out<=0;
   54595: out<=1;
   54596: out<=1;
   54597: out<=1;
   54598: out<=1;
   54599: out<=1;
   54600: out<=0;
   54601: out<=0;
   54602: out<=1;
   54603: out<=1;
   54604: out<=0;
   54605: out<=1;
   54606: out<=0;
   54607: out<=1;
   54608: out<=1;
   54609: out<=0;
   54610: out<=0;
   54611: out<=1;
   54612: out<=1;
   54613: out<=1;
   54614: out<=1;
   54615: out<=1;
   54616: out<=0;
   54617: out<=0;
   54618: out<=1;
   54619: out<=1;
   54620: out<=0;
   54621: out<=1;
   54622: out<=0;
   54623: out<=1;
   54624: out<=1;
   54625: out<=0;
   54626: out<=0;
   54627: out<=1;
   54628: out<=1;
   54629: out<=1;
   54630: out<=1;
   54631: out<=1;
   54632: out<=0;
   54633: out<=0;
   54634: out<=1;
   54635: out<=1;
   54636: out<=0;
   54637: out<=1;
   54638: out<=0;
   54639: out<=1;
   54640: out<=1;
   54641: out<=0;
   54642: out<=0;
   54643: out<=1;
   54644: out<=1;
   54645: out<=1;
   54646: out<=1;
   54647: out<=1;
   54648: out<=0;
   54649: out<=0;
   54650: out<=1;
   54651: out<=1;
   54652: out<=0;
   54653: out<=1;
   54654: out<=0;
   54655: out<=1;
   54656: out<=0;
   54657: out<=1;
   54658: out<=1;
   54659: out<=0;
   54660: out<=0;
   54661: out<=0;
   54662: out<=0;
   54663: out<=0;
   54664: out<=1;
   54665: out<=1;
   54666: out<=0;
   54667: out<=0;
   54668: out<=1;
   54669: out<=0;
   54670: out<=1;
   54671: out<=0;
   54672: out<=0;
   54673: out<=1;
   54674: out<=1;
   54675: out<=0;
   54676: out<=0;
   54677: out<=0;
   54678: out<=0;
   54679: out<=0;
   54680: out<=1;
   54681: out<=1;
   54682: out<=0;
   54683: out<=0;
   54684: out<=1;
   54685: out<=0;
   54686: out<=1;
   54687: out<=0;
   54688: out<=1;
   54689: out<=0;
   54690: out<=0;
   54691: out<=1;
   54692: out<=1;
   54693: out<=1;
   54694: out<=1;
   54695: out<=1;
   54696: out<=0;
   54697: out<=0;
   54698: out<=1;
   54699: out<=1;
   54700: out<=0;
   54701: out<=1;
   54702: out<=0;
   54703: out<=1;
   54704: out<=1;
   54705: out<=0;
   54706: out<=0;
   54707: out<=1;
   54708: out<=1;
   54709: out<=1;
   54710: out<=1;
   54711: out<=1;
   54712: out<=0;
   54713: out<=0;
   54714: out<=1;
   54715: out<=1;
   54716: out<=0;
   54717: out<=1;
   54718: out<=0;
   54719: out<=1;
   54720: out<=0;
   54721: out<=1;
   54722: out<=1;
   54723: out<=0;
   54724: out<=0;
   54725: out<=0;
   54726: out<=0;
   54727: out<=0;
   54728: out<=1;
   54729: out<=1;
   54730: out<=0;
   54731: out<=0;
   54732: out<=1;
   54733: out<=0;
   54734: out<=1;
   54735: out<=0;
   54736: out<=1;
   54737: out<=0;
   54738: out<=0;
   54739: out<=1;
   54740: out<=1;
   54741: out<=1;
   54742: out<=1;
   54743: out<=1;
   54744: out<=0;
   54745: out<=0;
   54746: out<=1;
   54747: out<=1;
   54748: out<=0;
   54749: out<=1;
   54750: out<=0;
   54751: out<=1;
   54752: out<=0;
   54753: out<=1;
   54754: out<=1;
   54755: out<=0;
   54756: out<=0;
   54757: out<=0;
   54758: out<=0;
   54759: out<=0;
   54760: out<=1;
   54761: out<=1;
   54762: out<=0;
   54763: out<=0;
   54764: out<=1;
   54765: out<=0;
   54766: out<=1;
   54767: out<=0;
   54768: out<=1;
   54769: out<=0;
   54770: out<=0;
   54771: out<=1;
   54772: out<=1;
   54773: out<=1;
   54774: out<=1;
   54775: out<=1;
   54776: out<=0;
   54777: out<=0;
   54778: out<=1;
   54779: out<=1;
   54780: out<=0;
   54781: out<=1;
   54782: out<=0;
   54783: out<=1;
   54784: out<=1;
   54785: out<=0;
   54786: out<=1;
   54787: out<=0;
   54788: out<=1;
   54789: out<=1;
   54790: out<=0;
   54791: out<=0;
   54792: out<=1;
   54793: out<=1;
   54794: out<=1;
   54795: out<=1;
   54796: out<=1;
   54797: out<=0;
   54798: out<=0;
   54799: out<=1;
   54800: out<=0;
   54801: out<=1;
   54802: out<=0;
   54803: out<=1;
   54804: out<=0;
   54805: out<=0;
   54806: out<=1;
   54807: out<=1;
   54808: out<=0;
   54809: out<=0;
   54810: out<=0;
   54811: out<=0;
   54812: out<=0;
   54813: out<=1;
   54814: out<=1;
   54815: out<=0;
   54816: out<=1;
   54817: out<=0;
   54818: out<=1;
   54819: out<=0;
   54820: out<=1;
   54821: out<=1;
   54822: out<=0;
   54823: out<=0;
   54824: out<=1;
   54825: out<=1;
   54826: out<=1;
   54827: out<=1;
   54828: out<=1;
   54829: out<=0;
   54830: out<=0;
   54831: out<=1;
   54832: out<=0;
   54833: out<=1;
   54834: out<=0;
   54835: out<=1;
   54836: out<=0;
   54837: out<=0;
   54838: out<=1;
   54839: out<=1;
   54840: out<=0;
   54841: out<=0;
   54842: out<=0;
   54843: out<=0;
   54844: out<=0;
   54845: out<=1;
   54846: out<=1;
   54847: out<=0;
   54848: out<=1;
   54849: out<=0;
   54850: out<=1;
   54851: out<=0;
   54852: out<=1;
   54853: out<=1;
   54854: out<=0;
   54855: out<=0;
   54856: out<=1;
   54857: out<=1;
   54858: out<=1;
   54859: out<=1;
   54860: out<=1;
   54861: out<=0;
   54862: out<=0;
   54863: out<=1;
   54864: out<=1;
   54865: out<=0;
   54866: out<=1;
   54867: out<=0;
   54868: out<=1;
   54869: out<=1;
   54870: out<=0;
   54871: out<=0;
   54872: out<=1;
   54873: out<=1;
   54874: out<=1;
   54875: out<=1;
   54876: out<=1;
   54877: out<=0;
   54878: out<=0;
   54879: out<=1;
   54880: out<=0;
   54881: out<=1;
   54882: out<=0;
   54883: out<=1;
   54884: out<=0;
   54885: out<=0;
   54886: out<=1;
   54887: out<=1;
   54888: out<=0;
   54889: out<=0;
   54890: out<=0;
   54891: out<=0;
   54892: out<=0;
   54893: out<=1;
   54894: out<=1;
   54895: out<=0;
   54896: out<=0;
   54897: out<=1;
   54898: out<=0;
   54899: out<=1;
   54900: out<=0;
   54901: out<=0;
   54902: out<=1;
   54903: out<=1;
   54904: out<=0;
   54905: out<=0;
   54906: out<=0;
   54907: out<=0;
   54908: out<=0;
   54909: out<=1;
   54910: out<=1;
   54911: out<=0;
   54912: out<=0;
   54913: out<=1;
   54914: out<=0;
   54915: out<=1;
   54916: out<=0;
   54917: out<=0;
   54918: out<=1;
   54919: out<=1;
   54920: out<=0;
   54921: out<=0;
   54922: out<=0;
   54923: out<=0;
   54924: out<=0;
   54925: out<=1;
   54926: out<=1;
   54927: out<=0;
   54928: out<=0;
   54929: out<=1;
   54930: out<=0;
   54931: out<=1;
   54932: out<=0;
   54933: out<=0;
   54934: out<=1;
   54935: out<=1;
   54936: out<=0;
   54937: out<=0;
   54938: out<=0;
   54939: out<=0;
   54940: out<=0;
   54941: out<=1;
   54942: out<=1;
   54943: out<=0;
   54944: out<=0;
   54945: out<=1;
   54946: out<=0;
   54947: out<=1;
   54948: out<=0;
   54949: out<=0;
   54950: out<=1;
   54951: out<=1;
   54952: out<=0;
   54953: out<=0;
   54954: out<=0;
   54955: out<=0;
   54956: out<=0;
   54957: out<=1;
   54958: out<=1;
   54959: out<=0;
   54960: out<=0;
   54961: out<=1;
   54962: out<=0;
   54963: out<=1;
   54964: out<=0;
   54965: out<=0;
   54966: out<=1;
   54967: out<=1;
   54968: out<=0;
   54969: out<=0;
   54970: out<=0;
   54971: out<=0;
   54972: out<=0;
   54973: out<=1;
   54974: out<=1;
   54975: out<=0;
   54976: out<=0;
   54977: out<=1;
   54978: out<=0;
   54979: out<=1;
   54980: out<=0;
   54981: out<=0;
   54982: out<=1;
   54983: out<=1;
   54984: out<=0;
   54985: out<=0;
   54986: out<=0;
   54987: out<=0;
   54988: out<=0;
   54989: out<=1;
   54990: out<=1;
   54991: out<=0;
   54992: out<=1;
   54993: out<=0;
   54994: out<=1;
   54995: out<=0;
   54996: out<=1;
   54997: out<=1;
   54998: out<=0;
   54999: out<=0;
   55000: out<=1;
   55001: out<=1;
   55002: out<=1;
   55003: out<=1;
   55004: out<=1;
   55005: out<=0;
   55006: out<=0;
   55007: out<=1;
   55008: out<=1;
   55009: out<=0;
   55010: out<=1;
   55011: out<=0;
   55012: out<=1;
   55013: out<=1;
   55014: out<=0;
   55015: out<=0;
   55016: out<=1;
   55017: out<=1;
   55018: out<=1;
   55019: out<=1;
   55020: out<=1;
   55021: out<=0;
   55022: out<=0;
   55023: out<=1;
   55024: out<=0;
   55025: out<=1;
   55026: out<=0;
   55027: out<=1;
   55028: out<=0;
   55029: out<=0;
   55030: out<=1;
   55031: out<=1;
   55032: out<=0;
   55033: out<=0;
   55034: out<=0;
   55035: out<=0;
   55036: out<=0;
   55037: out<=1;
   55038: out<=1;
   55039: out<=0;
   55040: out<=0;
   55041: out<=0;
   55042: out<=1;
   55043: out<=1;
   55044: out<=1;
   55045: out<=0;
   55046: out<=1;
   55047: out<=0;
   55048: out<=1;
   55049: out<=0;
   55050: out<=0;
   55051: out<=1;
   55052: out<=0;
   55053: out<=0;
   55054: out<=0;
   55055: out<=0;
   55056: out<=0;
   55057: out<=0;
   55058: out<=1;
   55059: out<=1;
   55060: out<=1;
   55061: out<=0;
   55062: out<=1;
   55063: out<=0;
   55064: out<=1;
   55065: out<=0;
   55066: out<=0;
   55067: out<=1;
   55068: out<=0;
   55069: out<=0;
   55070: out<=0;
   55071: out<=0;
   55072: out<=1;
   55073: out<=1;
   55074: out<=0;
   55075: out<=0;
   55076: out<=0;
   55077: out<=1;
   55078: out<=0;
   55079: out<=1;
   55080: out<=0;
   55081: out<=1;
   55082: out<=1;
   55083: out<=0;
   55084: out<=1;
   55085: out<=1;
   55086: out<=1;
   55087: out<=1;
   55088: out<=1;
   55089: out<=1;
   55090: out<=0;
   55091: out<=0;
   55092: out<=0;
   55093: out<=1;
   55094: out<=0;
   55095: out<=1;
   55096: out<=0;
   55097: out<=1;
   55098: out<=1;
   55099: out<=0;
   55100: out<=1;
   55101: out<=1;
   55102: out<=1;
   55103: out<=1;
   55104: out<=0;
   55105: out<=0;
   55106: out<=1;
   55107: out<=1;
   55108: out<=1;
   55109: out<=0;
   55110: out<=1;
   55111: out<=0;
   55112: out<=1;
   55113: out<=0;
   55114: out<=0;
   55115: out<=1;
   55116: out<=0;
   55117: out<=0;
   55118: out<=0;
   55119: out<=0;
   55120: out<=1;
   55121: out<=1;
   55122: out<=0;
   55123: out<=0;
   55124: out<=0;
   55125: out<=1;
   55126: out<=0;
   55127: out<=1;
   55128: out<=0;
   55129: out<=1;
   55130: out<=1;
   55131: out<=0;
   55132: out<=1;
   55133: out<=1;
   55134: out<=1;
   55135: out<=1;
   55136: out<=0;
   55137: out<=0;
   55138: out<=1;
   55139: out<=1;
   55140: out<=1;
   55141: out<=0;
   55142: out<=1;
   55143: out<=0;
   55144: out<=1;
   55145: out<=0;
   55146: out<=0;
   55147: out<=1;
   55148: out<=0;
   55149: out<=0;
   55150: out<=0;
   55151: out<=0;
   55152: out<=1;
   55153: out<=1;
   55154: out<=0;
   55155: out<=0;
   55156: out<=0;
   55157: out<=1;
   55158: out<=0;
   55159: out<=1;
   55160: out<=0;
   55161: out<=1;
   55162: out<=1;
   55163: out<=0;
   55164: out<=1;
   55165: out<=1;
   55166: out<=1;
   55167: out<=1;
   55168: out<=1;
   55169: out<=1;
   55170: out<=0;
   55171: out<=0;
   55172: out<=0;
   55173: out<=1;
   55174: out<=0;
   55175: out<=1;
   55176: out<=0;
   55177: out<=1;
   55178: out<=1;
   55179: out<=0;
   55180: out<=1;
   55181: out<=1;
   55182: out<=1;
   55183: out<=1;
   55184: out<=0;
   55185: out<=0;
   55186: out<=1;
   55187: out<=1;
   55188: out<=1;
   55189: out<=0;
   55190: out<=1;
   55191: out<=0;
   55192: out<=1;
   55193: out<=0;
   55194: out<=0;
   55195: out<=1;
   55196: out<=0;
   55197: out<=0;
   55198: out<=0;
   55199: out<=0;
   55200: out<=0;
   55201: out<=0;
   55202: out<=1;
   55203: out<=1;
   55204: out<=1;
   55205: out<=0;
   55206: out<=1;
   55207: out<=0;
   55208: out<=1;
   55209: out<=0;
   55210: out<=0;
   55211: out<=1;
   55212: out<=0;
   55213: out<=0;
   55214: out<=0;
   55215: out<=0;
   55216: out<=1;
   55217: out<=1;
   55218: out<=0;
   55219: out<=0;
   55220: out<=0;
   55221: out<=1;
   55222: out<=0;
   55223: out<=1;
   55224: out<=0;
   55225: out<=1;
   55226: out<=1;
   55227: out<=0;
   55228: out<=1;
   55229: out<=1;
   55230: out<=1;
   55231: out<=1;
   55232: out<=1;
   55233: out<=1;
   55234: out<=0;
   55235: out<=0;
   55236: out<=0;
   55237: out<=1;
   55238: out<=0;
   55239: out<=1;
   55240: out<=0;
   55241: out<=1;
   55242: out<=1;
   55243: out<=0;
   55244: out<=1;
   55245: out<=1;
   55246: out<=1;
   55247: out<=1;
   55248: out<=1;
   55249: out<=1;
   55250: out<=0;
   55251: out<=0;
   55252: out<=0;
   55253: out<=1;
   55254: out<=0;
   55255: out<=1;
   55256: out<=0;
   55257: out<=1;
   55258: out<=1;
   55259: out<=0;
   55260: out<=1;
   55261: out<=1;
   55262: out<=1;
   55263: out<=1;
   55264: out<=1;
   55265: out<=1;
   55266: out<=0;
   55267: out<=0;
   55268: out<=0;
   55269: out<=1;
   55270: out<=0;
   55271: out<=1;
   55272: out<=0;
   55273: out<=1;
   55274: out<=1;
   55275: out<=0;
   55276: out<=1;
   55277: out<=1;
   55278: out<=1;
   55279: out<=1;
   55280: out<=1;
   55281: out<=1;
   55282: out<=0;
   55283: out<=0;
   55284: out<=0;
   55285: out<=1;
   55286: out<=0;
   55287: out<=1;
   55288: out<=0;
   55289: out<=1;
   55290: out<=1;
   55291: out<=0;
   55292: out<=1;
   55293: out<=1;
   55294: out<=1;
   55295: out<=1;
   55296: out<=0;
   55297: out<=0;
   55298: out<=1;
   55299: out<=1;
   55300: out<=1;
   55301: out<=0;
   55302: out<=1;
   55303: out<=0;
   55304: out<=0;
   55305: out<=1;
   55306: out<=1;
   55307: out<=0;
   55308: out<=1;
   55309: out<=1;
   55310: out<=1;
   55311: out<=1;
   55312: out<=0;
   55313: out<=0;
   55314: out<=1;
   55315: out<=1;
   55316: out<=1;
   55317: out<=0;
   55318: out<=1;
   55319: out<=0;
   55320: out<=0;
   55321: out<=1;
   55322: out<=1;
   55323: out<=0;
   55324: out<=1;
   55325: out<=1;
   55326: out<=1;
   55327: out<=1;
   55328: out<=0;
   55329: out<=0;
   55330: out<=1;
   55331: out<=1;
   55332: out<=1;
   55333: out<=0;
   55334: out<=1;
   55335: out<=0;
   55336: out<=0;
   55337: out<=1;
   55338: out<=1;
   55339: out<=0;
   55340: out<=1;
   55341: out<=1;
   55342: out<=1;
   55343: out<=1;
   55344: out<=0;
   55345: out<=0;
   55346: out<=1;
   55347: out<=1;
   55348: out<=1;
   55349: out<=0;
   55350: out<=1;
   55351: out<=0;
   55352: out<=0;
   55353: out<=1;
   55354: out<=1;
   55355: out<=0;
   55356: out<=1;
   55357: out<=1;
   55358: out<=1;
   55359: out<=1;
   55360: out<=0;
   55361: out<=0;
   55362: out<=1;
   55363: out<=1;
   55364: out<=1;
   55365: out<=0;
   55366: out<=1;
   55367: out<=0;
   55368: out<=0;
   55369: out<=1;
   55370: out<=1;
   55371: out<=0;
   55372: out<=1;
   55373: out<=1;
   55374: out<=1;
   55375: out<=1;
   55376: out<=1;
   55377: out<=1;
   55378: out<=0;
   55379: out<=0;
   55380: out<=0;
   55381: out<=1;
   55382: out<=0;
   55383: out<=1;
   55384: out<=1;
   55385: out<=0;
   55386: out<=0;
   55387: out<=1;
   55388: out<=0;
   55389: out<=0;
   55390: out<=0;
   55391: out<=0;
   55392: out<=1;
   55393: out<=1;
   55394: out<=0;
   55395: out<=0;
   55396: out<=0;
   55397: out<=1;
   55398: out<=0;
   55399: out<=1;
   55400: out<=1;
   55401: out<=0;
   55402: out<=0;
   55403: out<=1;
   55404: out<=0;
   55405: out<=0;
   55406: out<=0;
   55407: out<=0;
   55408: out<=0;
   55409: out<=0;
   55410: out<=1;
   55411: out<=1;
   55412: out<=1;
   55413: out<=0;
   55414: out<=1;
   55415: out<=0;
   55416: out<=0;
   55417: out<=1;
   55418: out<=1;
   55419: out<=0;
   55420: out<=1;
   55421: out<=1;
   55422: out<=1;
   55423: out<=1;
   55424: out<=1;
   55425: out<=1;
   55426: out<=0;
   55427: out<=0;
   55428: out<=0;
   55429: out<=1;
   55430: out<=0;
   55431: out<=1;
   55432: out<=1;
   55433: out<=0;
   55434: out<=0;
   55435: out<=1;
   55436: out<=0;
   55437: out<=0;
   55438: out<=0;
   55439: out<=0;
   55440: out<=0;
   55441: out<=0;
   55442: out<=1;
   55443: out<=1;
   55444: out<=1;
   55445: out<=0;
   55446: out<=1;
   55447: out<=0;
   55448: out<=0;
   55449: out<=1;
   55450: out<=1;
   55451: out<=0;
   55452: out<=1;
   55453: out<=1;
   55454: out<=1;
   55455: out<=1;
   55456: out<=1;
   55457: out<=1;
   55458: out<=0;
   55459: out<=0;
   55460: out<=0;
   55461: out<=1;
   55462: out<=0;
   55463: out<=1;
   55464: out<=1;
   55465: out<=0;
   55466: out<=0;
   55467: out<=1;
   55468: out<=0;
   55469: out<=0;
   55470: out<=0;
   55471: out<=0;
   55472: out<=0;
   55473: out<=0;
   55474: out<=1;
   55475: out<=1;
   55476: out<=1;
   55477: out<=0;
   55478: out<=1;
   55479: out<=0;
   55480: out<=0;
   55481: out<=1;
   55482: out<=1;
   55483: out<=0;
   55484: out<=1;
   55485: out<=1;
   55486: out<=1;
   55487: out<=1;
   55488: out<=1;
   55489: out<=1;
   55490: out<=0;
   55491: out<=0;
   55492: out<=0;
   55493: out<=1;
   55494: out<=0;
   55495: out<=1;
   55496: out<=1;
   55497: out<=0;
   55498: out<=0;
   55499: out<=1;
   55500: out<=0;
   55501: out<=0;
   55502: out<=0;
   55503: out<=0;
   55504: out<=1;
   55505: out<=1;
   55506: out<=0;
   55507: out<=0;
   55508: out<=0;
   55509: out<=1;
   55510: out<=0;
   55511: out<=1;
   55512: out<=1;
   55513: out<=0;
   55514: out<=0;
   55515: out<=1;
   55516: out<=0;
   55517: out<=0;
   55518: out<=0;
   55519: out<=0;
   55520: out<=0;
   55521: out<=0;
   55522: out<=1;
   55523: out<=1;
   55524: out<=1;
   55525: out<=0;
   55526: out<=1;
   55527: out<=0;
   55528: out<=0;
   55529: out<=1;
   55530: out<=1;
   55531: out<=0;
   55532: out<=1;
   55533: out<=1;
   55534: out<=1;
   55535: out<=1;
   55536: out<=0;
   55537: out<=0;
   55538: out<=1;
   55539: out<=1;
   55540: out<=1;
   55541: out<=0;
   55542: out<=1;
   55543: out<=0;
   55544: out<=0;
   55545: out<=1;
   55546: out<=1;
   55547: out<=0;
   55548: out<=1;
   55549: out<=1;
   55550: out<=1;
   55551: out<=1;
   55552: out<=1;
   55553: out<=0;
   55554: out<=1;
   55555: out<=0;
   55556: out<=1;
   55557: out<=1;
   55558: out<=0;
   55559: out<=0;
   55560: out<=0;
   55561: out<=0;
   55562: out<=0;
   55563: out<=0;
   55564: out<=0;
   55565: out<=1;
   55566: out<=1;
   55567: out<=0;
   55568: out<=0;
   55569: out<=1;
   55570: out<=0;
   55571: out<=1;
   55572: out<=0;
   55573: out<=0;
   55574: out<=1;
   55575: out<=1;
   55576: out<=1;
   55577: out<=1;
   55578: out<=1;
   55579: out<=1;
   55580: out<=1;
   55581: out<=0;
   55582: out<=0;
   55583: out<=1;
   55584: out<=0;
   55585: out<=1;
   55586: out<=0;
   55587: out<=1;
   55588: out<=0;
   55589: out<=0;
   55590: out<=1;
   55591: out<=1;
   55592: out<=1;
   55593: out<=1;
   55594: out<=1;
   55595: out<=1;
   55596: out<=1;
   55597: out<=0;
   55598: out<=0;
   55599: out<=1;
   55600: out<=1;
   55601: out<=0;
   55602: out<=1;
   55603: out<=0;
   55604: out<=1;
   55605: out<=1;
   55606: out<=0;
   55607: out<=0;
   55608: out<=0;
   55609: out<=0;
   55610: out<=0;
   55611: out<=0;
   55612: out<=0;
   55613: out<=1;
   55614: out<=1;
   55615: out<=0;
   55616: out<=1;
   55617: out<=0;
   55618: out<=1;
   55619: out<=0;
   55620: out<=1;
   55621: out<=1;
   55622: out<=0;
   55623: out<=0;
   55624: out<=0;
   55625: out<=0;
   55626: out<=0;
   55627: out<=0;
   55628: out<=0;
   55629: out<=1;
   55630: out<=1;
   55631: out<=0;
   55632: out<=1;
   55633: out<=0;
   55634: out<=1;
   55635: out<=0;
   55636: out<=1;
   55637: out<=1;
   55638: out<=0;
   55639: out<=0;
   55640: out<=0;
   55641: out<=0;
   55642: out<=0;
   55643: out<=0;
   55644: out<=0;
   55645: out<=1;
   55646: out<=1;
   55647: out<=0;
   55648: out<=1;
   55649: out<=0;
   55650: out<=1;
   55651: out<=0;
   55652: out<=1;
   55653: out<=1;
   55654: out<=0;
   55655: out<=0;
   55656: out<=0;
   55657: out<=0;
   55658: out<=0;
   55659: out<=0;
   55660: out<=0;
   55661: out<=1;
   55662: out<=1;
   55663: out<=0;
   55664: out<=1;
   55665: out<=0;
   55666: out<=1;
   55667: out<=0;
   55668: out<=1;
   55669: out<=1;
   55670: out<=0;
   55671: out<=0;
   55672: out<=0;
   55673: out<=0;
   55674: out<=0;
   55675: out<=0;
   55676: out<=0;
   55677: out<=1;
   55678: out<=1;
   55679: out<=0;
   55680: out<=0;
   55681: out<=1;
   55682: out<=0;
   55683: out<=1;
   55684: out<=0;
   55685: out<=0;
   55686: out<=1;
   55687: out<=1;
   55688: out<=1;
   55689: out<=1;
   55690: out<=1;
   55691: out<=1;
   55692: out<=1;
   55693: out<=0;
   55694: out<=0;
   55695: out<=1;
   55696: out<=0;
   55697: out<=1;
   55698: out<=0;
   55699: out<=1;
   55700: out<=0;
   55701: out<=0;
   55702: out<=1;
   55703: out<=1;
   55704: out<=1;
   55705: out<=1;
   55706: out<=1;
   55707: out<=1;
   55708: out<=1;
   55709: out<=0;
   55710: out<=0;
   55711: out<=1;
   55712: out<=1;
   55713: out<=0;
   55714: out<=1;
   55715: out<=0;
   55716: out<=1;
   55717: out<=1;
   55718: out<=0;
   55719: out<=0;
   55720: out<=0;
   55721: out<=0;
   55722: out<=0;
   55723: out<=0;
   55724: out<=0;
   55725: out<=1;
   55726: out<=1;
   55727: out<=0;
   55728: out<=1;
   55729: out<=0;
   55730: out<=1;
   55731: out<=0;
   55732: out<=1;
   55733: out<=1;
   55734: out<=0;
   55735: out<=0;
   55736: out<=0;
   55737: out<=0;
   55738: out<=0;
   55739: out<=0;
   55740: out<=0;
   55741: out<=1;
   55742: out<=1;
   55743: out<=0;
   55744: out<=0;
   55745: out<=1;
   55746: out<=0;
   55747: out<=1;
   55748: out<=0;
   55749: out<=0;
   55750: out<=1;
   55751: out<=1;
   55752: out<=1;
   55753: out<=1;
   55754: out<=1;
   55755: out<=1;
   55756: out<=1;
   55757: out<=0;
   55758: out<=0;
   55759: out<=1;
   55760: out<=1;
   55761: out<=0;
   55762: out<=1;
   55763: out<=0;
   55764: out<=1;
   55765: out<=1;
   55766: out<=0;
   55767: out<=0;
   55768: out<=0;
   55769: out<=0;
   55770: out<=0;
   55771: out<=0;
   55772: out<=0;
   55773: out<=1;
   55774: out<=1;
   55775: out<=0;
   55776: out<=0;
   55777: out<=1;
   55778: out<=0;
   55779: out<=1;
   55780: out<=0;
   55781: out<=0;
   55782: out<=1;
   55783: out<=1;
   55784: out<=1;
   55785: out<=1;
   55786: out<=1;
   55787: out<=1;
   55788: out<=1;
   55789: out<=0;
   55790: out<=0;
   55791: out<=1;
   55792: out<=1;
   55793: out<=0;
   55794: out<=1;
   55795: out<=0;
   55796: out<=1;
   55797: out<=1;
   55798: out<=0;
   55799: out<=0;
   55800: out<=0;
   55801: out<=0;
   55802: out<=0;
   55803: out<=0;
   55804: out<=0;
   55805: out<=1;
   55806: out<=1;
   55807: out<=0;
   55808: out<=0;
   55809: out<=1;
   55810: out<=1;
   55811: out<=0;
   55812: out<=0;
   55813: out<=0;
   55814: out<=0;
   55815: out<=0;
   55816: out<=0;
   55817: out<=0;
   55818: out<=1;
   55819: out<=1;
   55820: out<=0;
   55821: out<=1;
   55822: out<=0;
   55823: out<=1;
   55824: out<=1;
   55825: out<=0;
   55826: out<=0;
   55827: out<=1;
   55828: out<=1;
   55829: out<=1;
   55830: out<=1;
   55831: out<=1;
   55832: out<=1;
   55833: out<=1;
   55834: out<=0;
   55835: out<=0;
   55836: out<=1;
   55837: out<=0;
   55838: out<=1;
   55839: out<=0;
   55840: out<=0;
   55841: out<=1;
   55842: out<=1;
   55843: out<=0;
   55844: out<=0;
   55845: out<=0;
   55846: out<=0;
   55847: out<=0;
   55848: out<=0;
   55849: out<=0;
   55850: out<=1;
   55851: out<=1;
   55852: out<=0;
   55853: out<=1;
   55854: out<=0;
   55855: out<=1;
   55856: out<=1;
   55857: out<=0;
   55858: out<=0;
   55859: out<=1;
   55860: out<=1;
   55861: out<=1;
   55862: out<=1;
   55863: out<=1;
   55864: out<=1;
   55865: out<=1;
   55866: out<=0;
   55867: out<=0;
   55868: out<=1;
   55869: out<=0;
   55870: out<=1;
   55871: out<=0;
   55872: out<=0;
   55873: out<=1;
   55874: out<=1;
   55875: out<=0;
   55876: out<=0;
   55877: out<=0;
   55878: out<=0;
   55879: out<=0;
   55880: out<=0;
   55881: out<=0;
   55882: out<=1;
   55883: out<=1;
   55884: out<=0;
   55885: out<=1;
   55886: out<=0;
   55887: out<=1;
   55888: out<=0;
   55889: out<=1;
   55890: out<=1;
   55891: out<=0;
   55892: out<=0;
   55893: out<=0;
   55894: out<=0;
   55895: out<=0;
   55896: out<=0;
   55897: out<=0;
   55898: out<=1;
   55899: out<=1;
   55900: out<=0;
   55901: out<=1;
   55902: out<=0;
   55903: out<=1;
   55904: out<=1;
   55905: out<=0;
   55906: out<=0;
   55907: out<=1;
   55908: out<=1;
   55909: out<=1;
   55910: out<=1;
   55911: out<=1;
   55912: out<=1;
   55913: out<=1;
   55914: out<=0;
   55915: out<=0;
   55916: out<=1;
   55917: out<=0;
   55918: out<=1;
   55919: out<=0;
   55920: out<=1;
   55921: out<=0;
   55922: out<=0;
   55923: out<=1;
   55924: out<=1;
   55925: out<=1;
   55926: out<=1;
   55927: out<=1;
   55928: out<=1;
   55929: out<=1;
   55930: out<=0;
   55931: out<=0;
   55932: out<=1;
   55933: out<=0;
   55934: out<=1;
   55935: out<=0;
   55936: out<=1;
   55937: out<=0;
   55938: out<=0;
   55939: out<=1;
   55940: out<=1;
   55941: out<=1;
   55942: out<=1;
   55943: out<=1;
   55944: out<=1;
   55945: out<=1;
   55946: out<=0;
   55947: out<=0;
   55948: out<=1;
   55949: out<=0;
   55950: out<=1;
   55951: out<=0;
   55952: out<=1;
   55953: out<=0;
   55954: out<=0;
   55955: out<=1;
   55956: out<=1;
   55957: out<=1;
   55958: out<=1;
   55959: out<=1;
   55960: out<=1;
   55961: out<=1;
   55962: out<=0;
   55963: out<=0;
   55964: out<=1;
   55965: out<=0;
   55966: out<=1;
   55967: out<=0;
   55968: out<=1;
   55969: out<=0;
   55970: out<=0;
   55971: out<=1;
   55972: out<=1;
   55973: out<=1;
   55974: out<=1;
   55975: out<=1;
   55976: out<=1;
   55977: out<=1;
   55978: out<=0;
   55979: out<=0;
   55980: out<=1;
   55981: out<=0;
   55982: out<=1;
   55983: out<=0;
   55984: out<=1;
   55985: out<=0;
   55986: out<=0;
   55987: out<=1;
   55988: out<=1;
   55989: out<=1;
   55990: out<=1;
   55991: out<=1;
   55992: out<=1;
   55993: out<=1;
   55994: out<=0;
   55995: out<=0;
   55996: out<=1;
   55997: out<=0;
   55998: out<=1;
   55999: out<=0;
   56000: out<=1;
   56001: out<=0;
   56002: out<=0;
   56003: out<=1;
   56004: out<=1;
   56005: out<=1;
   56006: out<=1;
   56007: out<=1;
   56008: out<=1;
   56009: out<=1;
   56010: out<=0;
   56011: out<=0;
   56012: out<=1;
   56013: out<=0;
   56014: out<=1;
   56015: out<=0;
   56016: out<=0;
   56017: out<=1;
   56018: out<=1;
   56019: out<=0;
   56020: out<=0;
   56021: out<=0;
   56022: out<=0;
   56023: out<=0;
   56024: out<=0;
   56025: out<=0;
   56026: out<=1;
   56027: out<=1;
   56028: out<=0;
   56029: out<=1;
   56030: out<=0;
   56031: out<=1;
   56032: out<=0;
   56033: out<=1;
   56034: out<=1;
   56035: out<=0;
   56036: out<=0;
   56037: out<=0;
   56038: out<=0;
   56039: out<=0;
   56040: out<=0;
   56041: out<=0;
   56042: out<=1;
   56043: out<=1;
   56044: out<=0;
   56045: out<=1;
   56046: out<=0;
   56047: out<=1;
   56048: out<=1;
   56049: out<=0;
   56050: out<=0;
   56051: out<=1;
   56052: out<=1;
   56053: out<=1;
   56054: out<=1;
   56055: out<=1;
   56056: out<=1;
   56057: out<=1;
   56058: out<=0;
   56059: out<=0;
   56060: out<=1;
   56061: out<=0;
   56062: out<=1;
   56063: out<=0;
   56064: out<=1;
   56065: out<=1;
   56066: out<=1;
   56067: out<=1;
   56068: out<=0;
   56069: out<=1;
   56070: out<=1;
   56071: out<=0;
   56072: out<=0;
   56073: out<=1;
   56074: out<=0;
   56075: out<=1;
   56076: out<=1;
   56077: out<=1;
   56078: out<=0;
   56079: out<=0;
   56080: out<=1;
   56081: out<=1;
   56082: out<=1;
   56083: out<=1;
   56084: out<=0;
   56085: out<=1;
   56086: out<=1;
   56087: out<=0;
   56088: out<=0;
   56089: out<=1;
   56090: out<=0;
   56091: out<=1;
   56092: out<=1;
   56093: out<=1;
   56094: out<=0;
   56095: out<=0;
   56096: out<=0;
   56097: out<=0;
   56098: out<=0;
   56099: out<=0;
   56100: out<=1;
   56101: out<=0;
   56102: out<=0;
   56103: out<=1;
   56104: out<=1;
   56105: out<=0;
   56106: out<=1;
   56107: out<=0;
   56108: out<=0;
   56109: out<=0;
   56110: out<=1;
   56111: out<=1;
   56112: out<=0;
   56113: out<=0;
   56114: out<=0;
   56115: out<=0;
   56116: out<=1;
   56117: out<=0;
   56118: out<=0;
   56119: out<=1;
   56120: out<=1;
   56121: out<=0;
   56122: out<=1;
   56123: out<=0;
   56124: out<=0;
   56125: out<=0;
   56126: out<=1;
   56127: out<=1;
   56128: out<=1;
   56129: out<=1;
   56130: out<=1;
   56131: out<=1;
   56132: out<=0;
   56133: out<=1;
   56134: out<=1;
   56135: out<=0;
   56136: out<=0;
   56137: out<=1;
   56138: out<=0;
   56139: out<=1;
   56140: out<=1;
   56141: out<=1;
   56142: out<=0;
   56143: out<=0;
   56144: out<=0;
   56145: out<=0;
   56146: out<=0;
   56147: out<=0;
   56148: out<=1;
   56149: out<=0;
   56150: out<=0;
   56151: out<=1;
   56152: out<=1;
   56153: out<=0;
   56154: out<=1;
   56155: out<=0;
   56156: out<=0;
   56157: out<=0;
   56158: out<=1;
   56159: out<=1;
   56160: out<=1;
   56161: out<=1;
   56162: out<=1;
   56163: out<=1;
   56164: out<=0;
   56165: out<=1;
   56166: out<=1;
   56167: out<=0;
   56168: out<=0;
   56169: out<=1;
   56170: out<=0;
   56171: out<=1;
   56172: out<=1;
   56173: out<=1;
   56174: out<=0;
   56175: out<=0;
   56176: out<=0;
   56177: out<=0;
   56178: out<=0;
   56179: out<=0;
   56180: out<=1;
   56181: out<=0;
   56182: out<=0;
   56183: out<=1;
   56184: out<=1;
   56185: out<=0;
   56186: out<=1;
   56187: out<=0;
   56188: out<=0;
   56189: out<=0;
   56190: out<=1;
   56191: out<=1;
   56192: out<=0;
   56193: out<=0;
   56194: out<=0;
   56195: out<=0;
   56196: out<=1;
   56197: out<=0;
   56198: out<=0;
   56199: out<=1;
   56200: out<=1;
   56201: out<=0;
   56202: out<=1;
   56203: out<=0;
   56204: out<=0;
   56205: out<=0;
   56206: out<=1;
   56207: out<=1;
   56208: out<=1;
   56209: out<=1;
   56210: out<=1;
   56211: out<=1;
   56212: out<=0;
   56213: out<=1;
   56214: out<=1;
   56215: out<=0;
   56216: out<=0;
   56217: out<=1;
   56218: out<=0;
   56219: out<=1;
   56220: out<=1;
   56221: out<=1;
   56222: out<=0;
   56223: out<=0;
   56224: out<=1;
   56225: out<=1;
   56226: out<=1;
   56227: out<=1;
   56228: out<=0;
   56229: out<=1;
   56230: out<=1;
   56231: out<=0;
   56232: out<=0;
   56233: out<=1;
   56234: out<=0;
   56235: out<=1;
   56236: out<=1;
   56237: out<=1;
   56238: out<=0;
   56239: out<=0;
   56240: out<=0;
   56241: out<=0;
   56242: out<=0;
   56243: out<=0;
   56244: out<=1;
   56245: out<=0;
   56246: out<=0;
   56247: out<=1;
   56248: out<=1;
   56249: out<=0;
   56250: out<=1;
   56251: out<=0;
   56252: out<=0;
   56253: out<=0;
   56254: out<=1;
   56255: out<=1;
   56256: out<=0;
   56257: out<=0;
   56258: out<=0;
   56259: out<=0;
   56260: out<=1;
   56261: out<=0;
   56262: out<=0;
   56263: out<=1;
   56264: out<=1;
   56265: out<=0;
   56266: out<=1;
   56267: out<=0;
   56268: out<=0;
   56269: out<=0;
   56270: out<=1;
   56271: out<=1;
   56272: out<=0;
   56273: out<=0;
   56274: out<=0;
   56275: out<=0;
   56276: out<=1;
   56277: out<=0;
   56278: out<=0;
   56279: out<=1;
   56280: out<=1;
   56281: out<=0;
   56282: out<=1;
   56283: out<=0;
   56284: out<=0;
   56285: out<=0;
   56286: out<=1;
   56287: out<=1;
   56288: out<=0;
   56289: out<=0;
   56290: out<=0;
   56291: out<=0;
   56292: out<=1;
   56293: out<=0;
   56294: out<=0;
   56295: out<=1;
   56296: out<=1;
   56297: out<=0;
   56298: out<=1;
   56299: out<=0;
   56300: out<=0;
   56301: out<=0;
   56302: out<=1;
   56303: out<=1;
   56304: out<=0;
   56305: out<=0;
   56306: out<=0;
   56307: out<=0;
   56308: out<=1;
   56309: out<=0;
   56310: out<=0;
   56311: out<=1;
   56312: out<=1;
   56313: out<=0;
   56314: out<=1;
   56315: out<=0;
   56316: out<=0;
   56317: out<=0;
   56318: out<=1;
   56319: out<=1;
   56320: out<=0;
   56321: out<=1;
   56322: out<=0;
   56323: out<=1;
   56324: out<=1;
   56325: out<=1;
   56326: out<=0;
   56327: out<=0;
   56328: out<=0;
   56329: out<=0;
   56330: out<=0;
   56331: out<=0;
   56332: out<=1;
   56333: out<=0;
   56334: out<=0;
   56335: out<=1;
   56336: out<=0;
   56337: out<=1;
   56338: out<=0;
   56339: out<=1;
   56340: out<=1;
   56341: out<=1;
   56342: out<=0;
   56343: out<=0;
   56344: out<=0;
   56345: out<=0;
   56346: out<=0;
   56347: out<=0;
   56348: out<=1;
   56349: out<=0;
   56350: out<=0;
   56351: out<=1;
   56352: out<=0;
   56353: out<=1;
   56354: out<=0;
   56355: out<=1;
   56356: out<=1;
   56357: out<=1;
   56358: out<=0;
   56359: out<=0;
   56360: out<=0;
   56361: out<=0;
   56362: out<=0;
   56363: out<=0;
   56364: out<=1;
   56365: out<=0;
   56366: out<=0;
   56367: out<=1;
   56368: out<=0;
   56369: out<=1;
   56370: out<=0;
   56371: out<=1;
   56372: out<=1;
   56373: out<=1;
   56374: out<=0;
   56375: out<=0;
   56376: out<=0;
   56377: out<=0;
   56378: out<=0;
   56379: out<=0;
   56380: out<=1;
   56381: out<=0;
   56382: out<=0;
   56383: out<=1;
   56384: out<=0;
   56385: out<=1;
   56386: out<=0;
   56387: out<=1;
   56388: out<=1;
   56389: out<=1;
   56390: out<=0;
   56391: out<=0;
   56392: out<=0;
   56393: out<=0;
   56394: out<=0;
   56395: out<=0;
   56396: out<=1;
   56397: out<=0;
   56398: out<=0;
   56399: out<=1;
   56400: out<=1;
   56401: out<=0;
   56402: out<=1;
   56403: out<=0;
   56404: out<=0;
   56405: out<=0;
   56406: out<=1;
   56407: out<=1;
   56408: out<=1;
   56409: out<=1;
   56410: out<=1;
   56411: out<=1;
   56412: out<=0;
   56413: out<=1;
   56414: out<=1;
   56415: out<=0;
   56416: out<=1;
   56417: out<=0;
   56418: out<=1;
   56419: out<=0;
   56420: out<=0;
   56421: out<=0;
   56422: out<=1;
   56423: out<=1;
   56424: out<=1;
   56425: out<=1;
   56426: out<=1;
   56427: out<=1;
   56428: out<=0;
   56429: out<=1;
   56430: out<=1;
   56431: out<=0;
   56432: out<=0;
   56433: out<=1;
   56434: out<=0;
   56435: out<=1;
   56436: out<=1;
   56437: out<=1;
   56438: out<=0;
   56439: out<=0;
   56440: out<=0;
   56441: out<=0;
   56442: out<=0;
   56443: out<=0;
   56444: out<=1;
   56445: out<=0;
   56446: out<=0;
   56447: out<=1;
   56448: out<=1;
   56449: out<=0;
   56450: out<=1;
   56451: out<=0;
   56452: out<=0;
   56453: out<=0;
   56454: out<=1;
   56455: out<=1;
   56456: out<=1;
   56457: out<=1;
   56458: out<=1;
   56459: out<=1;
   56460: out<=0;
   56461: out<=1;
   56462: out<=1;
   56463: out<=0;
   56464: out<=0;
   56465: out<=1;
   56466: out<=0;
   56467: out<=1;
   56468: out<=1;
   56469: out<=1;
   56470: out<=0;
   56471: out<=0;
   56472: out<=0;
   56473: out<=0;
   56474: out<=0;
   56475: out<=0;
   56476: out<=1;
   56477: out<=0;
   56478: out<=0;
   56479: out<=1;
   56480: out<=1;
   56481: out<=0;
   56482: out<=1;
   56483: out<=0;
   56484: out<=0;
   56485: out<=0;
   56486: out<=1;
   56487: out<=1;
   56488: out<=1;
   56489: out<=1;
   56490: out<=1;
   56491: out<=1;
   56492: out<=0;
   56493: out<=1;
   56494: out<=1;
   56495: out<=0;
   56496: out<=0;
   56497: out<=1;
   56498: out<=0;
   56499: out<=1;
   56500: out<=1;
   56501: out<=1;
   56502: out<=0;
   56503: out<=0;
   56504: out<=0;
   56505: out<=0;
   56506: out<=0;
   56507: out<=0;
   56508: out<=1;
   56509: out<=0;
   56510: out<=0;
   56511: out<=1;
   56512: out<=1;
   56513: out<=0;
   56514: out<=1;
   56515: out<=0;
   56516: out<=0;
   56517: out<=0;
   56518: out<=1;
   56519: out<=1;
   56520: out<=1;
   56521: out<=1;
   56522: out<=1;
   56523: out<=1;
   56524: out<=0;
   56525: out<=1;
   56526: out<=1;
   56527: out<=0;
   56528: out<=1;
   56529: out<=0;
   56530: out<=1;
   56531: out<=0;
   56532: out<=0;
   56533: out<=0;
   56534: out<=1;
   56535: out<=1;
   56536: out<=1;
   56537: out<=1;
   56538: out<=1;
   56539: out<=1;
   56540: out<=0;
   56541: out<=1;
   56542: out<=1;
   56543: out<=0;
   56544: out<=0;
   56545: out<=1;
   56546: out<=0;
   56547: out<=1;
   56548: out<=1;
   56549: out<=1;
   56550: out<=0;
   56551: out<=0;
   56552: out<=0;
   56553: out<=0;
   56554: out<=0;
   56555: out<=0;
   56556: out<=1;
   56557: out<=0;
   56558: out<=0;
   56559: out<=1;
   56560: out<=0;
   56561: out<=1;
   56562: out<=0;
   56563: out<=1;
   56564: out<=1;
   56565: out<=1;
   56566: out<=0;
   56567: out<=0;
   56568: out<=0;
   56569: out<=0;
   56570: out<=0;
   56571: out<=0;
   56572: out<=1;
   56573: out<=0;
   56574: out<=0;
   56575: out<=1;
   56576: out<=0;
   56577: out<=0;
   56578: out<=1;
   56579: out<=1;
   56580: out<=0;
   56581: out<=1;
   56582: out<=0;
   56583: out<=1;
   56584: out<=1;
   56585: out<=0;
   56586: out<=0;
   56587: out<=1;
   56588: out<=1;
   56589: out<=1;
   56590: out<=1;
   56591: out<=1;
   56592: out<=1;
   56593: out<=1;
   56594: out<=0;
   56595: out<=0;
   56596: out<=1;
   56597: out<=0;
   56598: out<=1;
   56599: out<=0;
   56600: out<=0;
   56601: out<=1;
   56602: out<=1;
   56603: out<=0;
   56604: out<=0;
   56605: out<=0;
   56606: out<=0;
   56607: out<=0;
   56608: out<=1;
   56609: out<=1;
   56610: out<=0;
   56611: out<=0;
   56612: out<=1;
   56613: out<=0;
   56614: out<=1;
   56615: out<=0;
   56616: out<=0;
   56617: out<=1;
   56618: out<=1;
   56619: out<=0;
   56620: out<=0;
   56621: out<=0;
   56622: out<=0;
   56623: out<=0;
   56624: out<=0;
   56625: out<=0;
   56626: out<=1;
   56627: out<=1;
   56628: out<=0;
   56629: out<=1;
   56630: out<=0;
   56631: out<=1;
   56632: out<=1;
   56633: out<=0;
   56634: out<=0;
   56635: out<=1;
   56636: out<=1;
   56637: out<=1;
   56638: out<=1;
   56639: out<=1;
   56640: out<=0;
   56641: out<=0;
   56642: out<=1;
   56643: out<=1;
   56644: out<=0;
   56645: out<=1;
   56646: out<=0;
   56647: out<=1;
   56648: out<=1;
   56649: out<=0;
   56650: out<=0;
   56651: out<=1;
   56652: out<=1;
   56653: out<=1;
   56654: out<=1;
   56655: out<=1;
   56656: out<=0;
   56657: out<=0;
   56658: out<=1;
   56659: out<=1;
   56660: out<=0;
   56661: out<=1;
   56662: out<=0;
   56663: out<=1;
   56664: out<=1;
   56665: out<=0;
   56666: out<=0;
   56667: out<=1;
   56668: out<=1;
   56669: out<=1;
   56670: out<=1;
   56671: out<=1;
   56672: out<=0;
   56673: out<=0;
   56674: out<=1;
   56675: out<=1;
   56676: out<=0;
   56677: out<=1;
   56678: out<=0;
   56679: out<=1;
   56680: out<=1;
   56681: out<=0;
   56682: out<=0;
   56683: out<=1;
   56684: out<=1;
   56685: out<=1;
   56686: out<=1;
   56687: out<=1;
   56688: out<=0;
   56689: out<=0;
   56690: out<=1;
   56691: out<=1;
   56692: out<=0;
   56693: out<=1;
   56694: out<=0;
   56695: out<=1;
   56696: out<=1;
   56697: out<=0;
   56698: out<=0;
   56699: out<=1;
   56700: out<=1;
   56701: out<=1;
   56702: out<=1;
   56703: out<=1;
   56704: out<=1;
   56705: out<=1;
   56706: out<=0;
   56707: out<=0;
   56708: out<=1;
   56709: out<=0;
   56710: out<=1;
   56711: out<=0;
   56712: out<=0;
   56713: out<=1;
   56714: out<=1;
   56715: out<=0;
   56716: out<=0;
   56717: out<=0;
   56718: out<=0;
   56719: out<=0;
   56720: out<=1;
   56721: out<=1;
   56722: out<=0;
   56723: out<=0;
   56724: out<=1;
   56725: out<=0;
   56726: out<=1;
   56727: out<=0;
   56728: out<=0;
   56729: out<=1;
   56730: out<=1;
   56731: out<=0;
   56732: out<=0;
   56733: out<=0;
   56734: out<=0;
   56735: out<=0;
   56736: out<=0;
   56737: out<=0;
   56738: out<=1;
   56739: out<=1;
   56740: out<=0;
   56741: out<=1;
   56742: out<=0;
   56743: out<=1;
   56744: out<=1;
   56745: out<=0;
   56746: out<=0;
   56747: out<=1;
   56748: out<=1;
   56749: out<=1;
   56750: out<=1;
   56751: out<=1;
   56752: out<=0;
   56753: out<=0;
   56754: out<=1;
   56755: out<=1;
   56756: out<=0;
   56757: out<=1;
   56758: out<=0;
   56759: out<=1;
   56760: out<=1;
   56761: out<=0;
   56762: out<=0;
   56763: out<=1;
   56764: out<=1;
   56765: out<=1;
   56766: out<=1;
   56767: out<=1;
   56768: out<=1;
   56769: out<=1;
   56770: out<=0;
   56771: out<=0;
   56772: out<=1;
   56773: out<=0;
   56774: out<=1;
   56775: out<=0;
   56776: out<=0;
   56777: out<=1;
   56778: out<=1;
   56779: out<=0;
   56780: out<=0;
   56781: out<=0;
   56782: out<=0;
   56783: out<=0;
   56784: out<=0;
   56785: out<=0;
   56786: out<=1;
   56787: out<=1;
   56788: out<=0;
   56789: out<=1;
   56790: out<=0;
   56791: out<=1;
   56792: out<=1;
   56793: out<=0;
   56794: out<=0;
   56795: out<=1;
   56796: out<=1;
   56797: out<=1;
   56798: out<=1;
   56799: out<=1;
   56800: out<=1;
   56801: out<=1;
   56802: out<=0;
   56803: out<=0;
   56804: out<=1;
   56805: out<=0;
   56806: out<=1;
   56807: out<=0;
   56808: out<=0;
   56809: out<=1;
   56810: out<=1;
   56811: out<=0;
   56812: out<=0;
   56813: out<=0;
   56814: out<=0;
   56815: out<=0;
   56816: out<=0;
   56817: out<=0;
   56818: out<=1;
   56819: out<=1;
   56820: out<=0;
   56821: out<=1;
   56822: out<=0;
   56823: out<=1;
   56824: out<=1;
   56825: out<=0;
   56826: out<=0;
   56827: out<=1;
   56828: out<=1;
   56829: out<=1;
   56830: out<=1;
   56831: out<=1;
   56832: out<=1;
   56833: out<=1;
   56834: out<=1;
   56835: out<=1;
   56836: out<=1;
   56837: out<=0;
   56838: out<=0;
   56839: out<=1;
   56840: out<=1;
   56841: out<=0;
   56842: out<=1;
   56843: out<=0;
   56844: out<=1;
   56845: out<=1;
   56846: out<=0;
   56847: out<=0;
   56848: out<=0;
   56849: out<=0;
   56850: out<=0;
   56851: out<=0;
   56852: out<=0;
   56853: out<=1;
   56854: out<=1;
   56855: out<=0;
   56856: out<=0;
   56857: out<=1;
   56858: out<=0;
   56859: out<=1;
   56860: out<=0;
   56861: out<=0;
   56862: out<=1;
   56863: out<=1;
   56864: out<=1;
   56865: out<=1;
   56866: out<=1;
   56867: out<=1;
   56868: out<=1;
   56869: out<=0;
   56870: out<=0;
   56871: out<=1;
   56872: out<=1;
   56873: out<=0;
   56874: out<=1;
   56875: out<=0;
   56876: out<=1;
   56877: out<=1;
   56878: out<=0;
   56879: out<=0;
   56880: out<=0;
   56881: out<=0;
   56882: out<=0;
   56883: out<=0;
   56884: out<=0;
   56885: out<=1;
   56886: out<=1;
   56887: out<=0;
   56888: out<=0;
   56889: out<=1;
   56890: out<=0;
   56891: out<=1;
   56892: out<=0;
   56893: out<=0;
   56894: out<=1;
   56895: out<=1;
   56896: out<=1;
   56897: out<=1;
   56898: out<=1;
   56899: out<=1;
   56900: out<=1;
   56901: out<=0;
   56902: out<=0;
   56903: out<=1;
   56904: out<=1;
   56905: out<=0;
   56906: out<=1;
   56907: out<=0;
   56908: out<=1;
   56909: out<=1;
   56910: out<=0;
   56911: out<=0;
   56912: out<=1;
   56913: out<=1;
   56914: out<=1;
   56915: out<=1;
   56916: out<=1;
   56917: out<=0;
   56918: out<=0;
   56919: out<=1;
   56920: out<=1;
   56921: out<=0;
   56922: out<=1;
   56923: out<=0;
   56924: out<=1;
   56925: out<=1;
   56926: out<=0;
   56927: out<=0;
   56928: out<=0;
   56929: out<=0;
   56930: out<=0;
   56931: out<=0;
   56932: out<=0;
   56933: out<=1;
   56934: out<=1;
   56935: out<=0;
   56936: out<=0;
   56937: out<=1;
   56938: out<=0;
   56939: out<=1;
   56940: out<=0;
   56941: out<=0;
   56942: out<=1;
   56943: out<=1;
   56944: out<=0;
   56945: out<=0;
   56946: out<=0;
   56947: out<=0;
   56948: out<=0;
   56949: out<=1;
   56950: out<=1;
   56951: out<=0;
   56952: out<=0;
   56953: out<=1;
   56954: out<=0;
   56955: out<=1;
   56956: out<=0;
   56957: out<=0;
   56958: out<=1;
   56959: out<=1;
   56960: out<=0;
   56961: out<=0;
   56962: out<=0;
   56963: out<=0;
   56964: out<=0;
   56965: out<=1;
   56966: out<=1;
   56967: out<=0;
   56968: out<=0;
   56969: out<=1;
   56970: out<=0;
   56971: out<=1;
   56972: out<=0;
   56973: out<=0;
   56974: out<=1;
   56975: out<=1;
   56976: out<=0;
   56977: out<=0;
   56978: out<=0;
   56979: out<=0;
   56980: out<=0;
   56981: out<=1;
   56982: out<=1;
   56983: out<=0;
   56984: out<=0;
   56985: out<=1;
   56986: out<=0;
   56987: out<=1;
   56988: out<=0;
   56989: out<=0;
   56990: out<=1;
   56991: out<=1;
   56992: out<=0;
   56993: out<=0;
   56994: out<=0;
   56995: out<=0;
   56996: out<=0;
   56997: out<=1;
   56998: out<=1;
   56999: out<=0;
   57000: out<=0;
   57001: out<=1;
   57002: out<=0;
   57003: out<=1;
   57004: out<=0;
   57005: out<=0;
   57006: out<=1;
   57007: out<=1;
   57008: out<=0;
   57009: out<=0;
   57010: out<=0;
   57011: out<=0;
   57012: out<=0;
   57013: out<=1;
   57014: out<=1;
   57015: out<=0;
   57016: out<=0;
   57017: out<=1;
   57018: out<=0;
   57019: out<=1;
   57020: out<=0;
   57021: out<=0;
   57022: out<=1;
   57023: out<=1;
   57024: out<=0;
   57025: out<=0;
   57026: out<=0;
   57027: out<=0;
   57028: out<=0;
   57029: out<=1;
   57030: out<=1;
   57031: out<=0;
   57032: out<=0;
   57033: out<=1;
   57034: out<=0;
   57035: out<=1;
   57036: out<=0;
   57037: out<=0;
   57038: out<=1;
   57039: out<=1;
   57040: out<=1;
   57041: out<=1;
   57042: out<=1;
   57043: out<=1;
   57044: out<=1;
   57045: out<=0;
   57046: out<=0;
   57047: out<=1;
   57048: out<=1;
   57049: out<=0;
   57050: out<=1;
   57051: out<=0;
   57052: out<=1;
   57053: out<=1;
   57054: out<=0;
   57055: out<=0;
   57056: out<=1;
   57057: out<=1;
   57058: out<=1;
   57059: out<=1;
   57060: out<=1;
   57061: out<=0;
   57062: out<=0;
   57063: out<=1;
   57064: out<=1;
   57065: out<=0;
   57066: out<=1;
   57067: out<=0;
   57068: out<=1;
   57069: out<=1;
   57070: out<=0;
   57071: out<=0;
   57072: out<=0;
   57073: out<=0;
   57074: out<=0;
   57075: out<=0;
   57076: out<=0;
   57077: out<=1;
   57078: out<=1;
   57079: out<=0;
   57080: out<=0;
   57081: out<=1;
   57082: out<=0;
   57083: out<=1;
   57084: out<=0;
   57085: out<=0;
   57086: out<=1;
   57087: out<=1;
   57088: out<=1;
   57089: out<=0;
   57090: out<=0;
   57091: out<=1;
   57092: out<=0;
   57093: out<=0;
   57094: out<=0;
   57095: out<=0;
   57096: out<=0;
   57097: out<=0;
   57098: out<=1;
   57099: out<=1;
   57100: out<=1;
   57101: out<=0;
   57102: out<=1;
   57103: out<=0;
   57104: out<=1;
   57105: out<=0;
   57106: out<=0;
   57107: out<=1;
   57108: out<=0;
   57109: out<=0;
   57110: out<=0;
   57111: out<=0;
   57112: out<=0;
   57113: out<=0;
   57114: out<=1;
   57115: out<=1;
   57116: out<=1;
   57117: out<=0;
   57118: out<=1;
   57119: out<=0;
   57120: out<=0;
   57121: out<=1;
   57122: out<=1;
   57123: out<=0;
   57124: out<=1;
   57125: out<=1;
   57126: out<=1;
   57127: out<=1;
   57128: out<=1;
   57129: out<=1;
   57130: out<=0;
   57131: out<=0;
   57132: out<=0;
   57133: out<=1;
   57134: out<=0;
   57135: out<=1;
   57136: out<=0;
   57137: out<=1;
   57138: out<=1;
   57139: out<=0;
   57140: out<=1;
   57141: out<=1;
   57142: out<=1;
   57143: out<=1;
   57144: out<=1;
   57145: out<=1;
   57146: out<=0;
   57147: out<=0;
   57148: out<=0;
   57149: out<=1;
   57150: out<=0;
   57151: out<=1;
   57152: out<=1;
   57153: out<=0;
   57154: out<=0;
   57155: out<=1;
   57156: out<=0;
   57157: out<=0;
   57158: out<=0;
   57159: out<=0;
   57160: out<=0;
   57161: out<=0;
   57162: out<=1;
   57163: out<=1;
   57164: out<=1;
   57165: out<=0;
   57166: out<=1;
   57167: out<=0;
   57168: out<=0;
   57169: out<=1;
   57170: out<=1;
   57171: out<=0;
   57172: out<=1;
   57173: out<=1;
   57174: out<=1;
   57175: out<=1;
   57176: out<=1;
   57177: out<=1;
   57178: out<=0;
   57179: out<=0;
   57180: out<=0;
   57181: out<=1;
   57182: out<=0;
   57183: out<=1;
   57184: out<=1;
   57185: out<=0;
   57186: out<=0;
   57187: out<=1;
   57188: out<=0;
   57189: out<=0;
   57190: out<=0;
   57191: out<=0;
   57192: out<=0;
   57193: out<=0;
   57194: out<=1;
   57195: out<=1;
   57196: out<=1;
   57197: out<=0;
   57198: out<=1;
   57199: out<=0;
   57200: out<=0;
   57201: out<=1;
   57202: out<=1;
   57203: out<=0;
   57204: out<=1;
   57205: out<=1;
   57206: out<=1;
   57207: out<=1;
   57208: out<=1;
   57209: out<=1;
   57210: out<=0;
   57211: out<=0;
   57212: out<=0;
   57213: out<=1;
   57214: out<=0;
   57215: out<=1;
   57216: out<=0;
   57217: out<=1;
   57218: out<=1;
   57219: out<=0;
   57220: out<=1;
   57221: out<=1;
   57222: out<=1;
   57223: out<=1;
   57224: out<=1;
   57225: out<=1;
   57226: out<=0;
   57227: out<=0;
   57228: out<=0;
   57229: out<=1;
   57230: out<=0;
   57231: out<=1;
   57232: out<=1;
   57233: out<=0;
   57234: out<=0;
   57235: out<=1;
   57236: out<=0;
   57237: out<=0;
   57238: out<=0;
   57239: out<=0;
   57240: out<=0;
   57241: out<=0;
   57242: out<=1;
   57243: out<=1;
   57244: out<=1;
   57245: out<=0;
   57246: out<=1;
   57247: out<=0;
   57248: out<=1;
   57249: out<=0;
   57250: out<=0;
   57251: out<=1;
   57252: out<=0;
   57253: out<=0;
   57254: out<=0;
   57255: out<=0;
   57256: out<=0;
   57257: out<=0;
   57258: out<=1;
   57259: out<=1;
   57260: out<=1;
   57261: out<=0;
   57262: out<=1;
   57263: out<=0;
   57264: out<=0;
   57265: out<=1;
   57266: out<=1;
   57267: out<=0;
   57268: out<=1;
   57269: out<=1;
   57270: out<=1;
   57271: out<=1;
   57272: out<=1;
   57273: out<=1;
   57274: out<=0;
   57275: out<=0;
   57276: out<=0;
   57277: out<=1;
   57278: out<=0;
   57279: out<=1;
   57280: out<=0;
   57281: out<=1;
   57282: out<=1;
   57283: out<=0;
   57284: out<=1;
   57285: out<=1;
   57286: out<=1;
   57287: out<=1;
   57288: out<=1;
   57289: out<=1;
   57290: out<=0;
   57291: out<=0;
   57292: out<=0;
   57293: out<=1;
   57294: out<=0;
   57295: out<=1;
   57296: out<=0;
   57297: out<=1;
   57298: out<=1;
   57299: out<=0;
   57300: out<=1;
   57301: out<=1;
   57302: out<=1;
   57303: out<=1;
   57304: out<=1;
   57305: out<=1;
   57306: out<=0;
   57307: out<=0;
   57308: out<=0;
   57309: out<=1;
   57310: out<=0;
   57311: out<=1;
   57312: out<=0;
   57313: out<=1;
   57314: out<=1;
   57315: out<=0;
   57316: out<=1;
   57317: out<=1;
   57318: out<=1;
   57319: out<=1;
   57320: out<=1;
   57321: out<=1;
   57322: out<=0;
   57323: out<=0;
   57324: out<=0;
   57325: out<=1;
   57326: out<=0;
   57327: out<=1;
   57328: out<=0;
   57329: out<=1;
   57330: out<=1;
   57331: out<=0;
   57332: out<=1;
   57333: out<=1;
   57334: out<=1;
   57335: out<=1;
   57336: out<=1;
   57337: out<=1;
   57338: out<=0;
   57339: out<=0;
   57340: out<=0;
   57341: out<=1;
   57342: out<=0;
   57343: out<=1;
   57344: out<=1;
   57345: out<=0;
   57346: out<=1;
   57347: out<=0;
   57348: out<=0;
   57349: out<=0;
   57350: out<=1;
   57351: out<=1;
   57352: out<=1;
   57353: out<=1;
   57354: out<=1;
   57355: out<=1;
   57356: out<=0;
   57357: out<=1;
   57358: out<=1;
   57359: out<=0;
   57360: out<=1;
   57361: out<=0;
   57362: out<=1;
   57363: out<=0;
   57364: out<=0;
   57365: out<=0;
   57366: out<=1;
   57367: out<=1;
   57368: out<=1;
   57369: out<=1;
   57370: out<=1;
   57371: out<=1;
   57372: out<=0;
   57373: out<=1;
   57374: out<=1;
   57375: out<=0;
   57376: out<=0;
   57377: out<=1;
   57378: out<=0;
   57379: out<=1;
   57380: out<=1;
   57381: out<=1;
   57382: out<=0;
   57383: out<=0;
   57384: out<=0;
   57385: out<=0;
   57386: out<=0;
   57387: out<=0;
   57388: out<=1;
   57389: out<=0;
   57390: out<=0;
   57391: out<=1;
   57392: out<=0;
   57393: out<=1;
   57394: out<=0;
   57395: out<=1;
   57396: out<=1;
   57397: out<=1;
   57398: out<=0;
   57399: out<=0;
   57400: out<=0;
   57401: out<=0;
   57402: out<=0;
   57403: out<=0;
   57404: out<=1;
   57405: out<=0;
   57406: out<=0;
   57407: out<=1;
   57408: out<=1;
   57409: out<=0;
   57410: out<=1;
   57411: out<=0;
   57412: out<=0;
   57413: out<=0;
   57414: out<=1;
   57415: out<=1;
   57416: out<=1;
   57417: out<=1;
   57418: out<=1;
   57419: out<=1;
   57420: out<=0;
   57421: out<=1;
   57422: out<=1;
   57423: out<=0;
   57424: out<=0;
   57425: out<=1;
   57426: out<=0;
   57427: out<=1;
   57428: out<=1;
   57429: out<=1;
   57430: out<=0;
   57431: out<=0;
   57432: out<=0;
   57433: out<=0;
   57434: out<=0;
   57435: out<=0;
   57436: out<=1;
   57437: out<=0;
   57438: out<=0;
   57439: out<=1;
   57440: out<=1;
   57441: out<=0;
   57442: out<=1;
   57443: out<=0;
   57444: out<=0;
   57445: out<=0;
   57446: out<=1;
   57447: out<=1;
   57448: out<=1;
   57449: out<=1;
   57450: out<=1;
   57451: out<=1;
   57452: out<=0;
   57453: out<=1;
   57454: out<=1;
   57455: out<=0;
   57456: out<=0;
   57457: out<=1;
   57458: out<=0;
   57459: out<=1;
   57460: out<=1;
   57461: out<=1;
   57462: out<=0;
   57463: out<=0;
   57464: out<=0;
   57465: out<=0;
   57466: out<=0;
   57467: out<=0;
   57468: out<=1;
   57469: out<=0;
   57470: out<=0;
   57471: out<=1;
   57472: out<=1;
   57473: out<=0;
   57474: out<=1;
   57475: out<=0;
   57476: out<=0;
   57477: out<=0;
   57478: out<=1;
   57479: out<=1;
   57480: out<=1;
   57481: out<=1;
   57482: out<=1;
   57483: out<=1;
   57484: out<=0;
   57485: out<=1;
   57486: out<=1;
   57487: out<=0;
   57488: out<=0;
   57489: out<=1;
   57490: out<=0;
   57491: out<=1;
   57492: out<=1;
   57493: out<=1;
   57494: out<=0;
   57495: out<=0;
   57496: out<=0;
   57497: out<=0;
   57498: out<=0;
   57499: out<=0;
   57500: out<=1;
   57501: out<=0;
   57502: out<=0;
   57503: out<=1;
   57504: out<=0;
   57505: out<=1;
   57506: out<=0;
   57507: out<=1;
   57508: out<=1;
   57509: out<=1;
   57510: out<=0;
   57511: out<=0;
   57512: out<=0;
   57513: out<=0;
   57514: out<=0;
   57515: out<=0;
   57516: out<=1;
   57517: out<=0;
   57518: out<=0;
   57519: out<=1;
   57520: out<=1;
   57521: out<=0;
   57522: out<=1;
   57523: out<=0;
   57524: out<=0;
   57525: out<=0;
   57526: out<=1;
   57527: out<=1;
   57528: out<=1;
   57529: out<=1;
   57530: out<=1;
   57531: out<=1;
   57532: out<=0;
   57533: out<=1;
   57534: out<=1;
   57535: out<=0;
   57536: out<=1;
   57537: out<=0;
   57538: out<=1;
   57539: out<=0;
   57540: out<=0;
   57541: out<=0;
   57542: out<=1;
   57543: out<=1;
   57544: out<=1;
   57545: out<=1;
   57546: out<=1;
   57547: out<=1;
   57548: out<=0;
   57549: out<=1;
   57550: out<=1;
   57551: out<=0;
   57552: out<=1;
   57553: out<=0;
   57554: out<=1;
   57555: out<=0;
   57556: out<=0;
   57557: out<=0;
   57558: out<=1;
   57559: out<=1;
   57560: out<=1;
   57561: out<=1;
   57562: out<=1;
   57563: out<=1;
   57564: out<=0;
   57565: out<=1;
   57566: out<=1;
   57567: out<=0;
   57568: out<=1;
   57569: out<=0;
   57570: out<=1;
   57571: out<=0;
   57572: out<=0;
   57573: out<=0;
   57574: out<=1;
   57575: out<=1;
   57576: out<=1;
   57577: out<=1;
   57578: out<=1;
   57579: out<=1;
   57580: out<=0;
   57581: out<=1;
   57582: out<=1;
   57583: out<=0;
   57584: out<=1;
   57585: out<=0;
   57586: out<=1;
   57587: out<=0;
   57588: out<=0;
   57589: out<=0;
   57590: out<=1;
   57591: out<=1;
   57592: out<=1;
   57593: out<=1;
   57594: out<=1;
   57595: out<=1;
   57596: out<=0;
   57597: out<=1;
   57598: out<=1;
   57599: out<=0;
   57600: out<=1;
   57601: out<=1;
   57602: out<=0;
   57603: out<=0;
   57604: out<=1;
   57605: out<=0;
   57606: out<=1;
   57607: out<=0;
   57608: out<=0;
   57609: out<=1;
   57610: out<=1;
   57611: out<=0;
   57612: out<=0;
   57613: out<=0;
   57614: out<=0;
   57615: out<=0;
   57616: out<=0;
   57617: out<=0;
   57618: out<=1;
   57619: out<=1;
   57620: out<=0;
   57621: out<=1;
   57622: out<=0;
   57623: out<=1;
   57624: out<=1;
   57625: out<=0;
   57626: out<=0;
   57627: out<=1;
   57628: out<=1;
   57629: out<=1;
   57630: out<=1;
   57631: out<=1;
   57632: out<=1;
   57633: out<=1;
   57634: out<=0;
   57635: out<=0;
   57636: out<=1;
   57637: out<=0;
   57638: out<=1;
   57639: out<=0;
   57640: out<=0;
   57641: out<=1;
   57642: out<=1;
   57643: out<=0;
   57644: out<=0;
   57645: out<=0;
   57646: out<=0;
   57647: out<=0;
   57648: out<=0;
   57649: out<=0;
   57650: out<=1;
   57651: out<=1;
   57652: out<=0;
   57653: out<=1;
   57654: out<=0;
   57655: out<=1;
   57656: out<=1;
   57657: out<=0;
   57658: out<=0;
   57659: out<=1;
   57660: out<=1;
   57661: out<=1;
   57662: out<=1;
   57663: out<=1;
   57664: out<=1;
   57665: out<=1;
   57666: out<=0;
   57667: out<=0;
   57668: out<=1;
   57669: out<=0;
   57670: out<=1;
   57671: out<=0;
   57672: out<=0;
   57673: out<=1;
   57674: out<=1;
   57675: out<=0;
   57676: out<=0;
   57677: out<=0;
   57678: out<=0;
   57679: out<=0;
   57680: out<=1;
   57681: out<=1;
   57682: out<=0;
   57683: out<=0;
   57684: out<=1;
   57685: out<=0;
   57686: out<=1;
   57687: out<=0;
   57688: out<=0;
   57689: out<=1;
   57690: out<=1;
   57691: out<=0;
   57692: out<=0;
   57693: out<=0;
   57694: out<=0;
   57695: out<=0;
   57696: out<=0;
   57697: out<=0;
   57698: out<=1;
   57699: out<=1;
   57700: out<=0;
   57701: out<=1;
   57702: out<=0;
   57703: out<=1;
   57704: out<=1;
   57705: out<=0;
   57706: out<=0;
   57707: out<=1;
   57708: out<=1;
   57709: out<=1;
   57710: out<=1;
   57711: out<=1;
   57712: out<=0;
   57713: out<=0;
   57714: out<=1;
   57715: out<=1;
   57716: out<=0;
   57717: out<=1;
   57718: out<=0;
   57719: out<=1;
   57720: out<=1;
   57721: out<=0;
   57722: out<=0;
   57723: out<=1;
   57724: out<=1;
   57725: out<=1;
   57726: out<=1;
   57727: out<=1;
   57728: out<=1;
   57729: out<=1;
   57730: out<=0;
   57731: out<=0;
   57732: out<=1;
   57733: out<=0;
   57734: out<=1;
   57735: out<=0;
   57736: out<=0;
   57737: out<=1;
   57738: out<=1;
   57739: out<=0;
   57740: out<=0;
   57741: out<=0;
   57742: out<=0;
   57743: out<=0;
   57744: out<=1;
   57745: out<=1;
   57746: out<=0;
   57747: out<=0;
   57748: out<=1;
   57749: out<=0;
   57750: out<=1;
   57751: out<=0;
   57752: out<=0;
   57753: out<=1;
   57754: out<=1;
   57755: out<=0;
   57756: out<=0;
   57757: out<=0;
   57758: out<=0;
   57759: out<=0;
   57760: out<=1;
   57761: out<=1;
   57762: out<=0;
   57763: out<=0;
   57764: out<=1;
   57765: out<=0;
   57766: out<=1;
   57767: out<=0;
   57768: out<=0;
   57769: out<=1;
   57770: out<=1;
   57771: out<=0;
   57772: out<=0;
   57773: out<=0;
   57774: out<=0;
   57775: out<=0;
   57776: out<=1;
   57777: out<=1;
   57778: out<=0;
   57779: out<=0;
   57780: out<=1;
   57781: out<=0;
   57782: out<=1;
   57783: out<=0;
   57784: out<=0;
   57785: out<=1;
   57786: out<=1;
   57787: out<=0;
   57788: out<=0;
   57789: out<=0;
   57790: out<=0;
   57791: out<=0;
   57792: out<=1;
   57793: out<=1;
   57794: out<=0;
   57795: out<=0;
   57796: out<=1;
   57797: out<=0;
   57798: out<=1;
   57799: out<=0;
   57800: out<=0;
   57801: out<=1;
   57802: out<=1;
   57803: out<=0;
   57804: out<=0;
   57805: out<=0;
   57806: out<=0;
   57807: out<=0;
   57808: out<=0;
   57809: out<=0;
   57810: out<=1;
   57811: out<=1;
   57812: out<=0;
   57813: out<=1;
   57814: out<=0;
   57815: out<=1;
   57816: out<=1;
   57817: out<=0;
   57818: out<=0;
   57819: out<=1;
   57820: out<=1;
   57821: out<=1;
   57822: out<=1;
   57823: out<=1;
   57824: out<=0;
   57825: out<=0;
   57826: out<=1;
   57827: out<=1;
   57828: out<=0;
   57829: out<=1;
   57830: out<=0;
   57831: out<=1;
   57832: out<=1;
   57833: out<=0;
   57834: out<=0;
   57835: out<=1;
   57836: out<=1;
   57837: out<=1;
   57838: out<=1;
   57839: out<=1;
   57840: out<=1;
   57841: out<=1;
   57842: out<=0;
   57843: out<=0;
   57844: out<=1;
   57845: out<=0;
   57846: out<=1;
   57847: out<=0;
   57848: out<=0;
   57849: out<=1;
   57850: out<=1;
   57851: out<=0;
   57852: out<=0;
   57853: out<=0;
   57854: out<=0;
   57855: out<=0;
   57856: out<=1;
   57857: out<=1;
   57858: out<=1;
   57859: out<=1;
   57860: out<=1;
   57861: out<=0;
   57862: out<=0;
   57863: out<=1;
   57864: out<=1;
   57865: out<=0;
   57866: out<=1;
   57867: out<=0;
   57868: out<=1;
   57869: out<=1;
   57870: out<=0;
   57871: out<=0;
   57872: out<=0;
   57873: out<=0;
   57874: out<=0;
   57875: out<=0;
   57876: out<=0;
   57877: out<=1;
   57878: out<=1;
   57879: out<=0;
   57880: out<=0;
   57881: out<=1;
   57882: out<=0;
   57883: out<=1;
   57884: out<=0;
   57885: out<=0;
   57886: out<=1;
   57887: out<=1;
   57888: out<=0;
   57889: out<=0;
   57890: out<=0;
   57891: out<=0;
   57892: out<=0;
   57893: out<=1;
   57894: out<=1;
   57895: out<=0;
   57896: out<=0;
   57897: out<=1;
   57898: out<=0;
   57899: out<=1;
   57900: out<=0;
   57901: out<=0;
   57902: out<=1;
   57903: out<=1;
   57904: out<=1;
   57905: out<=1;
   57906: out<=1;
   57907: out<=1;
   57908: out<=1;
   57909: out<=0;
   57910: out<=0;
   57911: out<=1;
   57912: out<=1;
   57913: out<=0;
   57914: out<=1;
   57915: out<=0;
   57916: out<=1;
   57917: out<=1;
   57918: out<=0;
   57919: out<=0;
   57920: out<=1;
   57921: out<=1;
   57922: out<=1;
   57923: out<=1;
   57924: out<=1;
   57925: out<=0;
   57926: out<=0;
   57927: out<=1;
   57928: out<=1;
   57929: out<=0;
   57930: out<=1;
   57931: out<=0;
   57932: out<=1;
   57933: out<=1;
   57934: out<=0;
   57935: out<=0;
   57936: out<=1;
   57937: out<=1;
   57938: out<=1;
   57939: out<=1;
   57940: out<=1;
   57941: out<=0;
   57942: out<=0;
   57943: out<=1;
   57944: out<=1;
   57945: out<=0;
   57946: out<=1;
   57947: out<=0;
   57948: out<=1;
   57949: out<=1;
   57950: out<=0;
   57951: out<=0;
   57952: out<=1;
   57953: out<=1;
   57954: out<=1;
   57955: out<=1;
   57956: out<=1;
   57957: out<=0;
   57958: out<=0;
   57959: out<=1;
   57960: out<=1;
   57961: out<=0;
   57962: out<=1;
   57963: out<=0;
   57964: out<=1;
   57965: out<=1;
   57966: out<=0;
   57967: out<=0;
   57968: out<=1;
   57969: out<=1;
   57970: out<=1;
   57971: out<=1;
   57972: out<=1;
   57973: out<=0;
   57974: out<=0;
   57975: out<=1;
   57976: out<=1;
   57977: out<=0;
   57978: out<=1;
   57979: out<=0;
   57980: out<=1;
   57981: out<=1;
   57982: out<=0;
   57983: out<=0;
   57984: out<=1;
   57985: out<=1;
   57986: out<=1;
   57987: out<=1;
   57988: out<=1;
   57989: out<=0;
   57990: out<=0;
   57991: out<=1;
   57992: out<=1;
   57993: out<=0;
   57994: out<=1;
   57995: out<=0;
   57996: out<=1;
   57997: out<=1;
   57998: out<=0;
   57999: out<=0;
   58000: out<=1;
   58001: out<=1;
   58002: out<=1;
   58003: out<=1;
   58004: out<=1;
   58005: out<=0;
   58006: out<=0;
   58007: out<=1;
   58008: out<=1;
   58009: out<=0;
   58010: out<=1;
   58011: out<=0;
   58012: out<=1;
   58013: out<=1;
   58014: out<=0;
   58015: out<=0;
   58016: out<=0;
   58017: out<=0;
   58018: out<=0;
   58019: out<=0;
   58020: out<=0;
   58021: out<=1;
   58022: out<=1;
   58023: out<=0;
   58024: out<=0;
   58025: out<=1;
   58026: out<=0;
   58027: out<=1;
   58028: out<=0;
   58029: out<=0;
   58030: out<=1;
   58031: out<=1;
   58032: out<=0;
   58033: out<=0;
   58034: out<=0;
   58035: out<=0;
   58036: out<=0;
   58037: out<=1;
   58038: out<=1;
   58039: out<=0;
   58040: out<=0;
   58041: out<=1;
   58042: out<=0;
   58043: out<=1;
   58044: out<=0;
   58045: out<=0;
   58046: out<=1;
   58047: out<=1;
   58048: out<=1;
   58049: out<=1;
   58050: out<=1;
   58051: out<=1;
   58052: out<=1;
   58053: out<=0;
   58054: out<=0;
   58055: out<=1;
   58056: out<=1;
   58057: out<=0;
   58058: out<=1;
   58059: out<=0;
   58060: out<=1;
   58061: out<=1;
   58062: out<=0;
   58063: out<=0;
   58064: out<=0;
   58065: out<=0;
   58066: out<=0;
   58067: out<=0;
   58068: out<=0;
   58069: out<=1;
   58070: out<=1;
   58071: out<=0;
   58072: out<=0;
   58073: out<=1;
   58074: out<=0;
   58075: out<=1;
   58076: out<=0;
   58077: out<=0;
   58078: out<=1;
   58079: out<=1;
   58080: out<=1;
   58081: out<=1;
   58082: out<=1;
   58083: out<=1;
   58084: out<=1;
   58085: out<=0;
   58086: out<=0;
   58087: out<=1;
   58088: out<=1;
   58089: out<=0;
   58090: out<=1;
   58091: out<=0;
   58092: out<=1;
   58093: out<=1;
   58094: out<=0;
   58095: out<=0;
   58096: out<=0;
   58097: out<=0;
   58098: out<=0;
   58099: out<=0;
   58100: out<=0;
   58101: out<=1;
   58102: out<=1;
   58103: out<=0;
   58104: out<=0;
   58105: out<=1;
   58106: out<=0;
   58107: out<=1;
   58108: out<=0;
   58109: out<=0;
   58110: out<=1;
   58111: out<=1;
   58112: out<=1;
   58113: out<=0;
   58114: out<=0;
   58115: out<=1;
   58116: out<=0;
   58117: out<=0;
   58118: out<=0;
   58119: out<=0;
   58120: out<=0;
   58121: out<=0;
   58122: out<=1;
   58123: out<=1;
   58124: out<=1;
   58125: out<=0;
   58126: out<=1;
   58127: out<=0;
   58128: out<=1;
   58129: out<=0;
   58130: out<=0;
   58131: out<=1;
   58132: out<=0;
   58133: out<=0;
   58134: out<=0;
   58135: out<=0;
   58136: out<=0;
   58137: out<=0;
   58138: out<=1;
   58139: out<=1;
   58140: out<=1;
   58141: out<=0;
   58142: out<=1;
   58143: out<=0;
   58144: out<=1;
   58145: out<=0;
   58146: out<=0;
   58147: out<=1;
   58148: out<=0;
   58149: out<=0;
   58150: out<=0;
   58151: out<=0;
   58152: out<=0;
   58153: out<=0;
   58154: out<=1;
   58155: out<=1;
   58156: out<=1;
   58157: out<=0;
   58158: out<=1;
   58159: out<=0;
   58160: out<=1;
   58161: out<=0;
   58162: out<=0;
   58163: out<=1;
   58164: out<=0;
   58165: out<=0;
   58166: out<=0;
   58167: out<=0;
   58168: out<=0;
   58169: out<=0;
   58170: out<=1;
   58171: out<=1;
   58172: out<=1;
   58173: out<=0;
   58174: out<=1;
   58175: out<=0;
   58176: out<=1;
   58177: out<=0;
   58178: out<=0;
   58179: out<=1;
   58180: out<=0;
   58181: out<=0;
   58182: out<=0;
   58183: out<=0;
   58184: out<=0;
   58185: out<=0;
   58186: out<=1;
   58187: out<=1;
   58188: out<=1;
   58189: out<=0;
   58190: out<=1;
   58191: out<=0;
   58192: out<=0;
   58193: out<=1;
   58194: out<=1;
   58195: out<=0;
   58196: out<=1;
   58197: out<=1;
   58198: out<=1;
   58199: out<=1;
   58200: out<=1;
   58201: out<=1;
   58202: out<=0;
   58203: out<=0;
   58204: out<=0;
   58205: out<=1;
   58206: out<=0;
   58207: out<=1;
   58208: out<=0;
   58209: out<=1;
   58210: out<=1;
   58211: out<=0;
   58212: out<=1;
   58213: out<=1;
   58214: out<=1;
   58215: out<=1;
   58216: out<=1;
   58217: out<=1;
   58218: out<=0;
   58219: out<=0;
   58220: out<=0;
   58221: out<=1;
   58222: out<=0;
   58223: out<=1;
   58224: out<=1;
   58225: out<=0;
   58226: out<=0;
   58227: out<=1;
   58228: out<=0;
   58229: out<=0;
   58230: out<=0;
   58231: out<=0;
   58232: out<=0;
   58233: out<=0;
   58234: out<=1;
   58235: out<=1;
   58236: out<=1;
   58237: out<=0;
   58238: out<=1;
   58239: out<=0;
   58240: out<=1;
   58241: out<=0;
   58242: out<=0;
   58243: out<=1;
   58244: out<=0;
   58245: out<=0;
   58246: out<=0;
   58247: out<=0;
   58248: out<=0;
   58249: out<=0;
   58250: out<=1;
   58251: out<=1;
   58252: out<=1;
   58253: out<=0;
   58254: out<=1;
   58255: out<=0;
   58256: out<=0;
   58257: out<=1;
   58258: out<=1;
   58259: out<=0;
   58260: out<=1;
   58261: out<=1;
   58262: out<=1;
   58263: out<=1;
   58264: out<=1;
   58265: out<=1;
   58266: out<=0;
   58267: out<=0;
   58268: out<=0;
   58269: out<=1;
   58270: out<=0;
   58271: out<=1;
   58272: out<=1;
   58273: out<=0;
   58274: out<=0;
   58275: out<=1;
   58276: out<=0;
   58277: out<=0;
   58278: out<=0;
   58279: out<=0;
   58280: out<=0;
   58281: out<=0;
   58282: out<=1;
   58283: out<=1;
   58284: out<=1;
   58285: out<=0;
   58286: out<=1;
   58287: out<=0;
   58288: out<=0;
   58289: out<=1;
   58290: out<=1;
   58291: out<=0;
   58292: out<=1;
   58293: out<=1;
   58294: out<=1;
   58295: out<=1;
   58296: out<=1;
   58297: out<=1;
   58298: out<=0;
   58299: out<=0;
   58300: out<=0;
   58301: out<=1;
   58302: out<=0;
   58303: out<=1;
   58304: out<=1;
   58305: out<=0;
   58306: out<=0;
   58307: out<=1;
   58308: out<=0;
   58309: out<=0;
   58310: out<=0;
   58311: out<=0;
   58312: out<=0;
   58313: out<=0;
   58314: out<=1;
   58315: out<=1;
   58316: out<=1;
   58317: out<=0;
   58318: out<=1;
   58319: out<=0;
   58320: out<=1;
   58321: out<=0;
   58322: out<=0;
   58323: out<=1;
   58324: out<=0;
   58325: out<=0;
   58326: out<=0;
   58327: out<=0;
   58328: out<=0;
   58329: out<=0;
   58330: out<=1;
   58331: out<=1;
   58332: out<=1;
   58333: out<=0;
   58334: out<=1;
   58335: out<=0;
   58336: out<=0;
   58337: out<=1;
   58338: out<=1;
   58339: out<=0;
   58340: out<=1;
   58341: out<=1;
   58342: out<=1;
   58343: out<=1;
   58344: out<=1;
   58345: out<=1;
   58346: out<=0;
   58347: out<=0;
   58348: out<=0;
   58349: out<=1;
   58350: out<=0;
   58351: out<=1;
   58352: out<=0;
   58353: out<=1;
   58354: out<=1;
   58355: out<=0;
   58356: out<=1;
   58357: out<=1;
   58358: out<=1;
   58359: out<=1;
   58360: out<=1;
   58361: out<=1;
   58362: out<=0;
   58363: out<=0;
   58364: out<=0;
   58365: out<=1;
   58366: out<=0;
   58367: out<=1;
   58368: out<=1;
   58369: out<=1;
   58370: out<=0;
   58371: out<=0;
   58372: out<=0;
   58373: out<=1;
   58374: out<=0;
   58375: out<=1;
   58376: out<=1;
   58377: out<=0;
   58378: out<=0;
   58379: out<=1;
   58380: out<=0;
   58381: out<=0;
   58382: out<=0;
   58383: out<=0;
   58384: out<=1;
   58385: out<=1;
   58386: out<=0;
   58387: out<=0;
   58388: out<=0;
   58389: out<=1;
   58390: out<=0;
   58391: out<=1;
   58392: out<=1;
   58393: out<=0;
   58394: out<=0;
   58395: out<=1;
   58396: out<=0;
   58397: out<=0;
   58398: out<=0;
   58399: out<=0;
   58400: out<=0;
   58401: out<=0;
   58402: out<=1;
   58403: out<=1;
   58404: out<=1;
   58405: out<=0;
   58406: out<=1;
   58407: out<=0;
   58408: out<=0;
   58409: out<=1;
   58410: out<=1;
   58411: out<=0;
   58412: out<=1;
   58413: out<=1;
   58414: out<=1;
   58415: out<=1;
   58416: out<=0;
   58417: out<=0;
   58418: out<=1;
   58419: out<=1;
   58420: out<=1;
   58421: out<=0;
   58422: out<=1;
   58423: out<=0;
   58424: out<=0;
   58425: out<=1;
   58426: out<=1;
   58427: out<=0;
   58428: out<=1;
   58429: out<=1;
   58430: out<=1;
   58431: out<=1;
   58432: out<=1;
   58433: out<=1;
   58434: out<=0;
   58435: out<=0;
   58436: out<=0;
   58437: out<=1;
   58438: out<=0;
   58439: out<=1;
   58440: out<=1;
   58441: out<=0;
   58442: out<=0;
   58443: out<=1;
   58444: out<=0;
   58445: out<=0;
   58446: out<=0;
   58447: out<=0;
   58448: out<=0;
   58449: out<=0;
   58450: out<=1;
   58451: out<=1;
   58452: out<=1;
   58453: out<=0;
   58454: out<=1;
   58455: out<=0;
   58456: out<=0;
   58457: out<=1;
   58458: out<=1;
   58459: out<=0;
   58460: out<=1;
   58461: out<=1;
   58462: out<=1;
   58463: out<=1;
   58464: out<=1;
   58465: out<=1;
   58466: out<=0;
   58467: out<=0;
   58468: out<=0;
   58469: out<=1;
   58470: out<=0;
   58471: out<=1;
   58472: out<=1;
   58473: out<=0;
   58474: out<=0;
   58475: out<=1;
   58476: out<=0;
   58477: out<=0;
   58478: out<=0;
   58479: out<=0;
   58480: out<=0;
   58481: out<=0;
   58482: out<=1;
   58483: out<=1;
   58484: out<=1;
   58485: out<=0;
   58486: out<=1;
   58487: out<=0;
   58488: out<=0;
   58489: out<=1;
   58490: out<=1;
   58491: out<=0;
   58492: out<=1;
   58493: out<=1;
   58494: out<=1;
   58495: out<=1;
   58496: out<=1;
   58497: out<=1;
   58498: out<=0;
   58499: out<=0;
   58500: out<=0;
   58501: out<=1;
   58502: out<=0;
   58503: out<=1;
   58504: out<=1;
   58505: out<=0;
   58506: out<=0;
   58507: out<=1;
   58508: out<=0;
   58509: out<=0;
   58510: out<=0;
   58511: out<=0;
   58512: out<=0;
   58513: out<=0;
   58514: out<=1;
   58515: out<=1;
   58516: out<=1;
   58517: out<=0;
   58518: out<=1;
   58519: out<=0;
   58520: out<=0;
   58521: out<=1;
   58522: out<=1;
   58523: out<=0;
   58524: out<=1;
   58525: out<=1;
   58526: out<=1;
   58527: out<=1;
   58528: out<=0;
   58529: out<=0;
   58530: out<=1;
   58531: out<=1;
   58532: out<=1;
   58533: out<=0;
   58534: out<=1;
   58535: out<=0;
   58536: out<=0;
   58537: out<=1;
   58538: out<=1;
   58539: out<=0;
   58540: out<=1;
   58541: out<=1;
   58542: out<=1;
   58543: out<=1;
   58544: out<=1;
   58545: out<=1;
   58546: out<=0;
   58547: out<=0;
   58548: out<=0;
   58549: out<=1;
   58550: out<=0;
   58551: out<=1;
   58552: out<=1;
   58553: out<=0;
   58554: out<=0;
   58555: out<=1;
   58556: out<=0;
   58557: out<=0;
   58558: out<=0;
   58559: out<=0;
   58560: out<=1;
   58561: out<=1;
   58562: out<=0;
   58563: out<=0;
   58564: out<=0;
   58565: out<=1;
   58566: out<=0;
   58567: out<=1;
   58568: out<=1;
   58569: out<=0;
   58570: out<=0;
   58571: out<=1;
   58572: out<=0;
   58573: out<=0;
   58574: out<=0;
   58575: out<=0;
   58576: out<=1;
   58577: out<=1;
   58578: out<=0;
   58579: out<=0;
   58580: out<=0;
   58581: out<=1;
   58582: out<=0;
   58583: out<=1;
   58584: out<=1;
   58585: out<=0;
   58586: out<=0;
   58587: out<=1;
   58588: out<=0;
   58589: out<=0;
   58590: out<=0;
   58591: out<=0;
   58592: out<=1;
   58593: out<=1;
   58594: out<=0;
   58595: out<=0;
   58596: out<=0;
   58597: out<=1;
   58598: out<=0;
   58599: out<=1;
   58600: out<=1;
   58601: out<=0;
   58602: out<=0;
   58603: out<=1;
   58604: out<=0;
   58605: out<=0;
   58606: out<=0;
   58607: out<=0;
   58608: out<=1;
   58609: out<=1;
   58610: out<=0;
   58611: out<=0;
   58612: out<=0;
   58613: out<=1;
   58614: out<=0;
   58615: out<=1;
   58616: out<=1;
   58617: out<=0;
   58618: out<=0;
   58619: out<=1;
   58620: out<=0;
   58621: out<=0;
   58622: out<=0;
   58623: out<=0;
   58624: out<=0;
   58625: out<=1;
   58626: out<=0;
   58627: out<=1;
   58628: out<=0;
   58629: out<=0;
   58630: out<=1;
   58631: out<=1;
   58632: out<=1;
   58633: out<=1;
   58634: out<=1;
   58635: out<=1;
   58636: out<=1;
   58637: out<=0;
   58638: out<=0;
   58639: out<=1;
   58640: out<=1;
   58641: out<=0;
   58642: out<=1;
   58643: out<=0;
   58644: out<=1;
   58645: out<=1;
   58646: out<=0;
   58647: out<=0;
   58648: out<=0;
   58649: out<=0;
   58650: out<=0;
   58651: out<=0;
   58652: out<=0;
   58653: out<=1;
   58654: out<=1;
   58655: out<=0;
   58656: out<=0;
   58657: out<=1;
   58658: out<=0;
   58659: out<=1;
   58660: out<=0;
   58661: out<=0;
   58662: out<=1;
   58663: out<=1;
   58664: out<=1;
   58665: out<=1;
   58666: out<=1;
   58667: out<=1;
   58668: out<=1;
   58669: out<=0;
   58670: out<=0;
   58671: out<=1;
   58672: out<=1;
   58673: out<=0;
   58674: out<=1;
   58675: out<=0;
   58676: out<=1;
   58677: out<=1;
   58678: out<=0;
   58679: out<=0;
   58680: out<=0;
   58681: out<=0;
   58682: out<=0;
   58683: out<=0;
   58684: out<=0;
   58685: out<=1;
   58686: out<=1;
   58687: out<=0;
   58688: out<=0;
   58689: out<=1;
   58690: out<=0;
   58691: out<=1;
   58692: out<=0;
   58693: out<=0;
   58694: out<=1;
   58695: out<=1;
   58696: out<=1;
   58697: out<=1;
   58698: out<=1;
   58699: out<=1;
   58700: out<=1;
   58701: out<=0;
   58702: out<=0;
   58703: out<=1;
   58704: out<=0;
   58705: out<=1;
   58706: out<=0;
   58707: out<=1;
   58708: out<=0;
   58709: out<=0;
   58710: out<=1;
   58711: out<=1;
   58712: out<=1;
   58713: out<=1;
   58714: out<=1;
   58715: out<=1;
   58716: out<=1;
   58717: out<=0;
   58718: out<=0;
   58719: out<=1;
   58720: out<=1;
   58721: out<=0;
   58722: out<=1;
   58723: out<=0;
   58724: out<=1;
   58725: out<=1;
   58726: out<=0;
   58727: out<=0;
   58728: out<=0;
   58729: out<=0;
   58730: out<=0;
   58731: out<=0;
   58732: out<=0;
   58733: out<=1;
   58734: out<=1;
   58735: out<=0;
   58736: out<=1;
   58737: out<=0;
   58738: out<=1;
   58739: out<=0;
   58740: out<=1;
   58741: out<=1;
   58742: out<=0;
   58743: out<=0;
   58744: out<=0;
   58745: out<=0;
   58746: out<=0;
   58747: out<=0;
   58748: out<=0;
   58749: out<=1;
   58750: out<=1;
   58751: out<=0;
   58752: out<=0;
   58753: out<=1;
   58754: out<=0;
   58755: out<=1;
   58756: out<=0;
   58757: out<=0;
   58758: out<=1;
   58759: out<=1;
   58760: out<=1;
   58761: out<=1;
   58762: out<=1;
   58763: out<=1;
   58764: out<=1;
   58765: out<=0;
   58766: out<=0;
   58767: out<=1;
   58768: out<=0;
   58769: out<=1;
   58770: out<=0;
   58771: out<=1;
   58772: out<=0;
   58773: out<=0;
   58774: out<=1;
   58775: out<=1;
   58776: out<=1;
   58777: out<=1;
   58778: out<=1;
   58779: out<=1;
   58780: out<=1;
   58781: out<=0;
   58782: out<=0;
   58783: out<=1;
   58784: out<=0;
   58785: out<=1;
   58786: out<=0;
   58787: out<=1;
   58788: out<=0;
   58789: out<=0;
   58790: out<=1;
   58791: out<=1;
   58792: out<=1;
   58793: out<=1;
   58794: out<=1;
   58795: out<=1;
   58796: out<=1;
   58797: out<=0;
   58798: out<=0;
   58799: out<=1;
   58800: out<=0;
   58801: out<=1;
   58802: out<=0;
   58803: out<=1;
   58804: out<=0;
   58805: out<=0;
   58806: out<=1;
   58807: out<=1;
   58808: out<=1;
   58809: out<=1;
   58810: out<=1;
   58811: out<=1;
   58812: out<=1;
   58813: out<=0;
   58814: out<=0;
   58815: out<=1;
   58816: out<=0;
   58817: out<=1;
   58818: out<=0;
   58819: out<=1;
   58820: out<=0;
   58821: out<=0;
   58822: out<=1;
   58823: out<=1;
   58824: out<=1;
   58825: out<=1;
   58826: out<=1;
   58827: out<=1;
   58828: out<=1;
   58829: out<=0;
   58830: out<=0;
   58831: out<=1;
   58832: out<=1;
   58833: out<=0;
   58834: out<=1;
   58835: out<=0;
   58836: out<=1;
   58837: out<=1;
   58838: out<=0;
   58839: out<=0;
   58840: out<=0;
   58841: out<=0;
   58842: out<=0;
   58843: out<=0;
   58844: out<=0;
   58845: out<=1;
   58846: out<=1;
   58847: out<=0;
   58848: out<=1;
   58849: out<=0;
   58850: out<=1;
   58851: out<=0;
   58852: out<=1;
   58853: out<=1;
   58854: out<=0;
   58855: out<=0;
   58856: out<=0;
   58857: out<=0;
   58858: out<=0;
   58859: out<=0;
   58860: out<=0;
   58861: out<=1;
   58862: out<=1;
   58863: out<=0;
   58864: out<=0;
   58865: out<=1;
   58866: out<=0;
   58867: out<=1;
   58868: out<=0;
   58869: out<=0;
   58870: out<=1;
   58871: out<=1;
   58872: out<=1;
   58873: out<=1;
   58874: out<=1;
   58875: out<=1;
   58876: out<=1;
   58877: out<=0;
   58878: out<=0;
   58879: out<=1;
   58880: out<=0;
   58881: out<=1;
   58882: out<=1;
   58883: out<=0;
   58884: out<=0;
   58885: out<=0;
   58886: out<=0;
   58887: out<=0;
   58888: out<=0;
   58889: out<=0;
   58890: out<=1;
   58891: out<=1;
   58892: out<=0;
   58893: out<=1;
   58894: out<=0;
   58895: out<=1;
   58896: out<=1;
   58897: out<=0;
   58898: out<=0;
   58899: out<=1;
   58900: out<=1;
   58901: out<=1;
   58902: out<=1;
   58903: out<=1;
   58904: out<=1;
   58905: out<=1;
   58906: out<=0;
   58907: out<=0;
   58908: out<=1;
   58909: out<=0;
   58910: out<=1;
   58911: out<=0;
   58912: out<=1;
   58913: out<=0;
   58914: out<=0;
   58915: out<=1;
   58916: out<=1;
   58917: out<=1;
   58918: out<=1;
   58919: out<=1;
   58920: out<=1;
   58921: out<=1;
   58922: out<=0;
   58923: out<=0;
   58924: out<=1;
   58925: out<=0;
   58926: out<=1;
   58927: out<=0;
   58928: out<=0;
   58929: out<=1;
   58930: out<=1;
   58931: out<=0;
   58932: out<=0;
   58933: out<=0;
   58934: out<=0;
   58935: out<=0;
   58936: out<=0;
   58937: out<=0;
   58938: out<=1;
   58939: out<=1;
   58940: out<=0;
   58941: out<=1;
   58942: out<=0;
   58943: out<=1;
   58944: out<=0;
   58945: out<=1;
   58946: out<=1;
   58947: out<=0;
   58948: out<=0;
   58949: out<=0;
   58950: out<=0;
   58951: out<=0;
   58952: out<=0;
   58953: out<=0;
   58954: out<=1;
   58955: out<=1;
   58956: out<=0;
   58957: out<=1;
   58958: out<=0;
   58959: out<=1;
   58960: out<=0;
   58961: out<=1;
   58962: out<=1;
   58963: out<=0;
   58964: out<=0;
   58965: out<=0;
   58966: out<=0;
   58967: out<=0;
   58968: out<=0;
   58969: out<=0;
   58970: out<=1;
   58971: out<=1;
   58972: out<=0;
   58973: out<=1;
   58974: out<=0;
   58975: out<=1;
   58976: out<=0;
   58977: out<=1;
   58978: out<=1;
   58979: out<=0;
   58980: out<=0;
   58981: out<=0;
   58982: out<=0;
   58983: out<=0;
   58984: out<=0;
   58985: out<=0;
   58986: out<=1;
   58987: out<=1;
   58988: out<=0;
   58989: out<=1;
   58990: out<=0;
   58991: out<=1;
   58992: out<=0;
   58993: out<=1;
   58994: out<=1;
   58995: out<=0;
   58996: out<=0;
   58997: out<=0;
   58998: out<=0;
   58999: out<=0;
   59000: out<=0;
   59001: out<=0;
   59002: out<=1;
   59003: out<=1;
   59004: out<=0;
   59005: out<=1;
   59006: out<=0;
   59007: out<=1;
   59008: out<=0;
   59009: out<=1;
   59010: out<=1;
   59011: out<=0;
   59012: out<=0;
   59013: out<=0;
   59014: out<=0;
   59015: out<=0;
   59016: out<=0;
   59017: out<=0;
   59018: out<=1;
   59019: out<=1;
   59020: out<=0;
   59021: out<=1;
   59022: out<=0;
   59023: out<=1;
   59024: out<=0;
   59025: out<=1;
   59026: out<=1;
   59027: out<=0;
   59028: out<=0;
   59029: out<=0;
   59030: out<=0;
   59031: out<=0;
   59032: out<=0;
   59033: out<=0;
   59034: out<=1;
   59035: out<=1;
   59036: out<=0;
   59037: out<=1;
   59038: out<=0;
   59039: out<=1;
   59040: out<=1;
   59041: out<=0;
   59042: out<=0;
   59043: out<=1;
   59044: out<=1;
   59045: out<=1;
   59046: out<=1;
   59047: out<=1;
   59048: out<=1;
   59049: out<=1;
   59050: out<=0;
   59051: out<=0;
   59052: out<=1;
   59053: out<=0;
   59054: out<=1;
   59055: out<=0;
   59056: out<=1;
   59057: out<=0;
   59058: out<=0;
   59059: out<=1;
   59060: out<=1;
   59061: out<=1;
   59062: out<=1;
   59063: out<=1;
   59064: out<=1;
   59065: out<=1;
   59066: out<=0;
   59067: out<=0;
   59068: out<=1;
   59069: out<=0;
   59070: out<=1;
   59071: out<=0;
   59072: out<=0;
   59073: out<=1;
   59074: out<=1;
   59075: out<=0;
   59076: out<=0;
   59077: out<=0;
   59078: out<=0;
   59079: out<=0;
   59080: out<=0;
   59081: out<=0;
   59082: out<=1;
   59083: out<=1;
   59084: out<=0;
   59085: out<=1;
   59086: out<=0;
   59087: out<=1;
   59088: out<=1;
   59089: out<=0;
   59090: out<=0;
   59091: out<=1;
   59092: out<=1;
   59093: out<=1;
   59094: out<=1;
   59095: out<=1;
   59096: out<=1;
   59097: out<=1;
   59098: out<=0;
   59099: out<=0;
   59100: out<=1;
   59101: out<=0;
   59102: out<=1;
   59103: out<=0;
   59104: out<=0;
   59105: out<=1;
   59106: out<=1;
   59107: out<=0;
   59108: out<=0;
   59109: out<=0;
   59110: out<=0;
   59111: out<=0;
   59112: out<=0;
   59113: out<=0;
   59114: out<=1;
   59115: out<=1;
   59116: out<=0;
   59117: out<=1;
   59118: out<=0;
   59119: out<=1;
   59120: out<=1;
   59121: out<=0;
   59122: out<=0;
   59123: out<=1;
   59124: out<=1;
   59125: out<=1;
   59126: out<=1;
   59127: out<=1;
   59128: out<=1;
   59129: out<=1;
   59130: out<=0;
   59131: out<=0;
   59132: out<=1;
   59133: out<=0;
   59134: out<=1;
   59135: out<=0;
   59136: out<=1;
   59137: out<=1;
   59138: out<=1;
   59139: out<=1;
   59140: out<=0;
   59141: out<=1;
   59142: out<=1;
   59143: out<=0;
   59144: out<=0;
   59145: out<=1;
   59146: out<=0;
   59147: out<=1;
   59148: out<=1;
   59149: out<=1;
   59150: out<=0;
   59151: out<=0;
   59152: out<=1;
   59153: out<=1;
   59154: out<=1;
   59155: out<=1;
   59156: out<=0;
   59157: out<=1;
   59158: out<=1;
   59159: out<=0;
   59160: out<=0;
   59161: out<=1;
   59162: out<=0;
   59163: out<=1;
   59164: out<=1;
   59165: out<=1;
   59166: out<=0;
   59167: out<=0;
   59168: out<=1;
   59169: out<=1;
   59170: out<=1;
   59171: out<=1;
   59172: out<=0;
   59173: out<=1;
   59174: out<=1;
   59175: out<=0;
   59176: out<=0;
   59177: out<=1;
   59178: out<=0;
   59179: out<=1;
   59180: out<=1;
   59181: out<=1;
   59182: out<=0;
   59183: out<=0;
   59184: out<=1;
   59185: out<=1;
   59186: out<=1;
   59187: out<=1;
   59188: out<=0;
   59189: out<=1;
   59190: out<=1;
   59191: out<=0;
   59192: out<=0;
   59193: out<=1;
   59194: out<=0;
   59195: out<=1;
   59196: out<=1;
   59197: out<=1;
   59198: out<=0;
   59199: out<=0;
   59200: out<=1;
   59201: out<=1;
   59202: out<=1;
   59203: out<=1;
   59204: out<=0;
   59205: out<=1;
   59206: out<=1;
   59207: out<=0;
   59208: out<=0;
   59209: out<=1;
   59210: out<=0;
   59211: out<=1;
   59212: out<=1;
   59213: out<=1;
   59214: out<=0;
   59215: out<=0;
   59216: out<=0;
   59217: out<=0;
   59218: out<=0;
   59219: out<=0;
   59220: out<=1;
   59221: out<=0;
   59222: out<=0;
   59223: out<=1;
   59224: out<=1;
   59225: out<=0;
   59226: out<=1;
   59227: out<=0;
   59228: out<=0;
   59229: out<=0;
   59230: out<=1;
   59231: out<=1;
   59232: out<=0;
   59233: out<=0;
   59234: out<=0;
   59235: out<=0;
   59236: out<=1;
   59237: out<=0;
   59238: out<=0;
   59239: out<=1;
   59240: out<=1;
   59241: out<=0;
   59242: out<=1;
   59243: out<=0;
   59244: out<=0;
   59245: out<=0;
   59246: out<=1;
   59247: out<=1;
   59248: out<=1;
   59249: out<=1;
   59250: out<=1;
   59251: out<=1;
   59252: out<=0;
   59253: out<=1;
   59254: out<=1;
   59255: out<=0;
   59256: out<=0;
   59257: out<=1;
   59258: out<=0;
   59259: out<=1;
   59260: out<=1;
   59261: out<=1;
   59262: out<=0;
   59263: out<=0;
   59264: out<=1;
   59265: out<=1;
   59266: out<=1;
   59267: out<=1;
   59268: out<=0;
   59269: out<=1;
   59270: out<=1;
   59271: out<=0;
   59272: out<=0;
   59273: out<=1;
   59274: out<=0;
   59275: out<=1;
   59276: out<=1;
   59277: out<=1;
   59278: out<=0;
   59279: out<=0;
   59280: out<=0;
   59281: out<=0;
   59282: out<=0;
   59283: out<=0;
   59284: out<=1;
   59285: out<=0;
   59286: out<=0;
   59287: out<=1;
   59288: out<=1;
   59289: out<=0;
   59290: out<=1;
   59291: out<=0;
   59292: out<=0;
   59293: out<=0;
   59294: out<=1;
   59295: out<=1;
   59296: out<=1;
   59297: out<=1;
   59298: out<=1;
   59299: out<=1;
   59300: out<=0;
   59301: out<=1;
   59302: out<=1;
   59303: out<=0;
   59304: out<=0;
   59305: out<=1;
   59306: out<=0;
   59307: out<=1;
   59308: out<=1;
   59309: out<=1;
   59310: out<=0;
   59311: out<=0;
   59312: out<=0;
   59313: out<=0;
   59314: out<=0;
   59315: out<=0;
   59316: out<=1;
   59317: out<=0;
   59318: out<=0;
   59319: out<=1;
   59320: out<=1;
   59321: out<=0;
   59322: out<=1;
   59323: out<=0;
   59324: out<=0;
   59325: out<=0;
   59326: out<=1;
   59327: out<=1;
   59328: out<=1;
   59329: out<=1;
   59330: out<=1;
   59331: out<=1;
   59332: out<=0;
   59333: out<=1;
   59334: out<=1;
   59335: out<=0;
   59336: out<=0;
   59337: out<=1;
   59338: out<=0;
   59339: out<=1;
   59340: out<=1;
   59341: out<=1;
   59342: out<=0;
   59343: out<=0;
   59344: out<=1;
   59345: out<=1;
   59346: out<=1;
   59347: out<=1;
   59348: out<=0;
   59349: out<=1;
   59350: out<=1;
   59351: out<=0;
   59352: out<=0;
   59353: out<=1;
   59354: out<=0;
   59355: out<=1;
   59356: out<=1;
   59357: out<=1;
   59358: out<=0;
   59359: out<=0;
   59360: out<=0;
   59361: out<=0;
   59362: out<=0;
   59363: out<=0;
   59364: out<=1;
   59365: out<=0;
   59366: out<=0;
   59367: out<=1;
   59368: out<=1;
   59369: out<=0;
   59370: out<=1;
   59371: out<=0;
   59372: out<=0;
   59373: out<=0;
   59374: out<=1;
   59375: out<=1;
   59376: out<=0;
   59377: out<=0;
   59378: out<=0;
   59379: out<=0;
   59380: out<=1;
   59381: out<=0;
   59382: out<=0;
   59383: out<=1;
   59384: out<=1;
   59385: out<=0;
   59386: out<=1;
   59387: out<=0;
   59388: out<=0;
   59389: out<=0;
   59390: out<=1;
   59391: out<=1;
   59392: out<=1;
   59393: out<=1;
   59394: out<=1;
   59395: out<=1;
   59396: out<=0;
   59397: out<=1;
   59398: out<=1;
   59399: out<=0;
   59400: out<=1;
   59401: out<=0;
   59402: out<=1;
   59403: out<=0;
   59404: out<=0;
   59405: out<=0;
   59406: out<=1;
   59407: out<=1;
   59408: out<=1;
   59409: out<=1;
   59410: out<=1;
   59411: out<=1;
   59412: out<=0;
   59413: out<=1;
   59414: out<=1;
   59415: out<=0;
   59416: out<=1;
   59417: out<=0;
   59418: out<=1;
   59419: out<=0;
   59420: out<=0;
   59421: out<=0;
   59422: out<=1;
   59423: out<=1;
   59424: out<=0;
   59425: out<=0;
   59426: out<=0;
   59427: out<=0;
   59428: out<=1;
   59429: out<=0;
   59430: out<=0;
   59431: out<=1;
   59432: out<=0;
   59433: out<=1;
   59434: out<=0;
   59435: out<=1;
   59436: out<=1;
   59437: out<=1;
   59438: out<=0;
   59439: out<=0;
   59440: out<=0;
   59441: out<=0;
   59442: out<=0;
   59443: out<=0;
   59444: out<=1;
   59445: out<=0;
   59446: out<=0;
   59447: out<=1;
   59448: out<=0;
   59449: out<=1;
   59450: out<=0;
   59451: out<=1;
   59452: out<=1;
   59453: out<=1;
   59454: out<=0;
   59455: out<=0;
   59456: out<=1;
   59457: out<=1;
   59458: out<=1;
   59459: out<=1;
   59460: out<=0;
   59461: out<=1;
   59462: out<=1;
   59463: out<=0;
   59464: out<=1;
   59465: out<=0;
   59466: out<=1;
   59467: out<=0;
   59468: out<=0;
   59469: out<=0;
   59470: out<=1;
   59471: out<=1;
   59472: out<=0;
   59473: out<=0;
   59474: out<=0;
   59475: out<=0;
   59476: out<=1;
   59477: out<=0;
   59478: out<=0;
   59479: out<=1;
   59480: out<=0;
   59481: out<=1;
   59482: out<=0;
   59483: out<=1;
   59484: out<=1;
   59485: out<=1;
   59486: out<=0;
   59487: out<=0;
   59488: out<=1;
   59489: out<=1;
   59490: out<=1;
   59491: out<=1;
   59492: out<=0;
   59493: out<=1;
   59494: out<=1;
   59495: out<=0;
   59496: out<=1;
   59497: out<=0;
   59498: out<=1;
   59499: out<=0;
   59500: out<=0;
   59501: out<=0;
   59502: out<=1;
   59503: out<=1;
   59504: out<=0;
   59505: out<=0;
   59506: out<=0;
   59507: out<=0;
   59508: out<=1;
   59509: out<=0;
   59510: out<=0;
   59511: out<=1;
   59512: out<=0;
   59513: out<=1;
   59514: out<=0;
   59515: out<=1;
   59516: out<=1;
   59517: out<=1;
   59518: out<=0;
   59519: out<=0;
   59520: out<=1;
   59521: out<=1;
   59522: out<=1;
   59523: out<=1;
   59524: out<=0;
   59525: out<=1;
   59526: out<=1;
   59527: out<=0;
   59528: out<=1;
   59529: out<=0;
   59530: out<=1;
   59531: out<=0;
   59532: out<=0;
   59533: out<=0;
   59534: out<=1;
   59535: out<=1;
   59536: out<=0;
   59537: out<=0;
   59538: out<=0;
   59539: out<=0;
   59540: out<=1;
   59541: out<=0;
   59542: out<=0;
   59543: out<=1;
   59544: out<=0;
   59545: out<=1;
   59546: out<=0;
   59547: out<=1;
   59548: out<=1;
   59549: out<=1;
   59550: out<=0;
   59551: out<=0;
   59552: out<=0;
   59553: out<=0;
   59554: out<=0;
   59555: out<=0;
   59556: out<=1;
   59557: out<=0;
   59558: out<=0;
   59559: out<=1;
   59560: out<=0;
   59561: out<=1;
   59562: out<=0;
   59563: out<=1;
   59564: out<=1;
   59565: out<=1;
   59566: out<=0;
   59567: out<=0;
   59568: out<=1;
   59569: out<=1;
   59570: out<=1;
   59571: out<=1;
   59572: out<=0;
   59573: out<=1;
   59574: out<=1;
   59575: out<=0;
   59576: out<=1;
   59577: out<=0;
   59578: out<=1;
   59579: out<=0;
   59580: out<=0;
   59581: out<=0;
   59582: out<=1;
   59583: out<=1;
   59584: out<=1;
   59585: out<=1;
   59586: out<=1;
   59587: out<=1;
   59588: out<=0;
   59589: out<=1;
   59590: out<=1;
   59591: out<=0;
   59592: out<=1;
   59593: out<=0;
   59594: out<=1;
   59595: out<=0;
   59596: out<=0;
   59597: out<=0;
   59598: out<=1;
   59599: out<=1;
   59600: out<=1;
   59601: out<=1;
   59602: out<=1;
   59603: out<=1;
   59604: out<=0;
   59605: out<=1;
   59606: out<=1;
   59607: out<=0;
   59608: out<=1;
   59609: out<=0;
   59610: out<=1;
   59611: out<=0;
   59612: out<=0;
   59613: out<=0;
   59614: out<=1;
   59615: out<=1;
   59616: out<=1;
   59617: out<=1;
   59618: out<=1;
   59619: out<=1;
   59620: out<=0;
   59621: out<=1;
   59622: out<=1;
   59623: out<=0;
   59624: out<=1;
   59625: out<=0;
   59626: out<=1;
   59627: out<=0;
   59628: out<=0;
   59629: out<=0;
   59630: out<=1;
   59631: out<=1;
   59632: out<=1;
   59633: out<=1;
   59634: out<=1;
   59635: out<=1;
   59636: out<=0;
   59637: out<=1;
   59638: out<=1;
   59639: out<=0;
   59640: out<=1;
   59641: out<=0;
   59642: out<=1;
   59643: out<=0;
   59644: out<=0;
   59645: out<=0;
   59646: out<=1;
   59647: out<=1;
   59648: out<=0;
   59649: out<=1;
   59650: out<=1;
   59651: out<=0;
   59652: out<=0;
   59653: out<=0;
   59654: out<=0;
   59655: out<=0;
   59656: out<=1;
   59657: out<=1;
   59658: out<=0;
   59659: out<=0;
   59660: out<=1;
   59661: out<=0;
   59662: out<=1;
   59663: out<=0;
   59664: out<=1;
   59665: out<=0;
   59666: out<=0;
   59667: out<=1;
   59668: out<=1;
   59669: out<=1;
   59670: out<=1;
   59671: out<=1;
   59672: out<=0;
   59673: out<=0;
   59674: out<=1;
   59675: out<=1;
   59676: out<=0;
   59677: out<=1;
   59678: out<=0;
   59679: out<=1;
   59680: out<=0;
   59681: out<=1;
   59682: out<=1;
   59683: out<=0;
   59684: out<=0;
   59685: out<=0;
   59686: out<=0;
   59687: out<=0;
   59688: out<=1;
   59689: out<=1;
   59690: out<=0;
   59691: out<=0;
   59692: out<=1;
   59693: out<=0;
   59694: out<=1;
   59695: out<=0;
   59696: out<=1;
   59697: out<=0;
   59698: out<=0;
   59699: out<=1;
   59700: out<=1;
   59701: out<=1;
   59702: out<=1;
   59703: out<=1;
   59704: out<=0;
   59705: out<=0;
   59706: out<=1;
   59707: out<=1;
   59708: out<=0;
   59709: out<=1;
   59710: out<=0;
   59711: out<=1;
   59712: out<=0;
   59713: out<=1;
   59714: out<=1;
   59715: out<=0;
   59716: out<=0;
   59717: out<=0;
   59718: out<=0;
   59719: out<=0;
   59720: out<=1;
   59721: out<=1;
   59722: out<=0;
   59723: out<=0;
   59724: out<=1;
   59725: out<=0;
   59726: out<=1;
   59727: out<=0;
   59728: out<=0;
   59729: out<=1;
   59730: out<=1;
   59731: out<=0;
   59732: out<=0;
   59733: out<=0;
   59734: out<=0;
   59735: out<=0;
   59736: out<=1;
   59737: out<=1;
   59738: out<=0;
   59739: out<=0;
   59740: out<=1;
   59741: out<=0;
   59742: out<=1;
   59743: out<=0;
   59744: out<=1;
   59745: out<=0;
   59746: out<=0;
   59747: out<=1;
   59748: out<=1;
   59749: out<=1;
   59750: out<=1;
   59751: out<=1;
   59752: out<=0;
   59753: out<=0;
   59754: out<=1;
   59755: out<=1;
   59756: out<=0;
   59757: out<=1;
   59758: out<=0;
   59759: out<=1;
   59760: out<=1;
   59761: out<=0;
   59762: out<=0;
   59763: out<=1;
   59764: out<=1;
   59765: out<=1;
   59766: out<=1;
   59767: out<=1;
   59768: out<=0;
   59769: out<=0;
   59770: out<=1;
   59771: out<=1;
   59772: out<=0;
   59773: out<=1;
   59774: out<=0;
   59775: out<=1;
   59776: out<=0;
   59777: out<=1;
   59778: out<=1;
   59779: out<=0;
   59780: out<=0;
   59781: out<=0;
   59782: out<=0;
   59783: out<=0;
   59784: out<=1;
   59785: out<=1;
   59786: out<=0;
   59787: out<=0;
   59788: out<=1;
   59789: out<=0;
   59790: out<=1;
   59791: out<=0;
   59792: out<=0;
   59793: out<=1;
   59794: out<=1;
   59795: out<=0;
   59796: out<=0;
   59797: out<=0;
   59798: out<=0;
   59799: out<=0;
   59800: out<=1;
   59801: out<=1;
   59802: out<=0;
   59803: out<=0;
   59804: out<=1;
   59805: out<=0;
   59806: out<=1;
   59807: out<=0;
   59808: out<=0;
   59809: out<=1;
   59810: out<=1;
   59811: out<=0;
   59812: out<=0;
   59813: out<=0;
   59814: out<=0;
   59815: out<=0;
   59816: out<=1;
   59817: out<=1;
   59818: out<=0;
   59819: out<=0;
   59820: out<=1;
   59821: out<=0;
   59822: out<=1;
   59823: out<=0;
   59824: out<=0;
   59825: out<=1;
   59826: out<=1;
   59827: out<=0;
   59828: out<=0;
   59829: out<=0;
   59830: out<=0;
   59831: out<=0;
   59832: out<=1;
   59833: out<=1;
   59834: out<=0;
   59835: out<=0;
   59836: out<=1;
   59837: out<=0;
   59838: out<=1;
   59839: out<=0;
   59840: out<=0;
   59841: out<=1;
   59842: out<=1;
   59843: out<=0;
   59844: out<=0;
   59845: out<=0;
   59846: out<=0;
   59847: out<=0;
   59848: out<=1;
   59849: out<=1;
   59850: out<=0;
   59851: out<=0;
   59852: out<=1;
   59853: out<=0;
   59854: out<=1;
   59855: out<=0;
   59856: out<=1;
   59857: out<=0;
   59858: out<=0;
   59859: out<=1;
   59860: out<=1;
   59861: out<=1;
   59862: out<=1;
   59863: out<=1;
   59864: out<=0;
   59865: out<=0;
   59866: out<=1;
   59867: out<=1;
   59868: out<=0;
   59869: out<=1;
   59870: out<=0;
   59871: out<=1;
   59872: out<=1;
   59873: out<=0;
   59874: out<=0;
   59875: out<=1;
   59876: out<=1;
   59877: out<=1;
   59878: out<=1;
   59879: out<=1;
   59880: out<=0;
   59881: out<=0;
   59882: out<=1;
   59883: out<=1;
   59884: out<=0;
   59885: out<=1;
   59886: out<=0;
   59887: out<=1;
   59888: out<=0;
   59889: out<=1;
   59890: out<=1;
   59891: out<=0;
   59892: out<=0;
   59893: out<=0;
   59894: out<=0;
   59895: out<=0;
   59896: out<=1;
   59897: out<=1;
   59898: out<=0;
   59899: out<=0;
   59900: out<=1;
   59901: out<=0;
   59902: out<=1;
   59903: out<=0;
   59904: out<=1;
   59905: out<=0;
   59906: out<=1;
   59907: out<=0;
   59908: out<=1;
   59909: out<=1;
   59910: out<=0;
   59911: out<=0;
   59912: out<=1;
   59913: out<=1;
   59914: out<=1;
   59915: out<=1;
   59916: out<=1;
   59917: out<=0;
   59918: out<=0;
   59919: out<=1;
   59920: out<=0;
   59921: out<=1;
   59922: out<=0;
   59923: out<=1;
   59924: out<=0;
   59925: out<=0;
   59926: out<=1;
   59927: out<=1;
   59928: out<=0;
   59929: out<=0;
   59930: out<=0;
   59931: out<=0;
   59932: out<=0;
   59933: out<=1;
   59934: out<=1;
   59935: out<=0;
   59936: out<=0;
   59937: out<=1;
   59938: out<=0;
   59939: out<=1;
   59940: out<=0;
   59941: out<=0;
   59942: out<=1;
   59943: out<=1;
   59944: out<=0;
   59945: out<=0;
   59946: out<=0;
   59947: out<=0;
   59948: out<=0;
   59949: out<=1;
   59950: out<=1;
   59951: out<=0;
   59952: out<=1;
   59953: out<=0;
   59954: out<=1;
   59955: out<=0;
   59956: out<=1;
   59957: out<=1;
   59958: out<=0;
   59959: out<=0;
   59960: out<=1;
   59961: out<=1;
   59962: out<=1;
   59963: out<=1;
   59964: out<=1;
   59965: out<=0;
   59966: out<=0;
   59967: out<=1;
   59968: out<=1;
   59969: out<=0;
   59970: out<=1;
   59971: out<=0;
   59972: out<=1;
   59973: out<=1;
   59974: out<=0;
   59975: out<=0;
   59976: out<=1;
   59977: out<=1;
   59978: out<=1;
   59979: out<=1;
   59980: out<=1;
   59981: out<=0;
   59982: out<=0;
   59983: out<=1;
   59984: out<=1;
   59985: out<=0;
   59986: out<=1;
   59987: out<=0;
   59988: out<=1;
   59989: out<=1;
   59990: out<=0;
   59991: out<=0;
   59992: out<=1;
   59993: out<=1;
   59994: out<=1;
   59995: out<=1;
   59996: out<=1;
   59997: out<=0;
   59998: out<=0;
   59999: out<=1;
   60000: out<=1;
   60001: out<=0;
   60002: out<=1;
   60003: out<=0;
   60004: out<=1;
   60005: out<=1;
   60006: out<=0;
   60007: out<=0;
   60008: out<=1;
   60009: out<=1;
   60010: out<=1;
   60011: out<=1;
   60012: out<=1;
   60013: out<=0;
   60014: out<=0;
   60015: out<=1;
   60016: out<=1;
   60017: out<=0;
   60018: out<=1;
   60019: out<=0;
   60020: out<=1;
   60021: out<=1;
   60022: out<=0;
   60023: out<=0;
   60024: out<=1;
   60025: out<=1;
   60026: out<=1;
   60027: out<=1;
   60028: out<=1;
   60029: out<=0;
   60030: out<=0;
   60031: out<=1;
   60032: out<=1;
   60033: out<=0;
   60034: out<=1;
   60035: out<=0;
   60036: out<=1;
   60037: out<=1;
   60038: out<=0;
   60039: out<=0;
   60040: out<=1;
   60041: out<=1;
   60042: out<=1;
   60043: out<=1;
   60044: out<=1;
   60045: out<=0;
   60046: out<=0;
   60047: out<=1;
   60048: out<=1;
   60049: out<=0;
   60050: out<=1;
   60051: out<=0;
   60052: out<=1;
   60053: out<=1;
   60054: out<=0;
   60055: out<=0;
   60056: out<=1;
   60057: out<=1;
   60058: out<=1;
   60059: out<=1;
   60060: out<=1;
   60061: out<=0;
   60062: out<=0;
   60063: out<=1;
   60064: out<=0;
   60065: out<=1;
   60066: out<=0;
   60067: out<=1;
   60068: out<=0;
   60069: out<=0;
   60070: out<=1;
   60071: out<=1;
   60072: out<=0;
   60073: out<=0;
   60074: out<=0;
   60075: out<=0;
   60076: out<=0;
   60077: out<=1;
   60078: out<=1;
   60079: out<=0;
   60080: out<=0;
   60081: out<=1;
   60082: out<=0;
   60083: out<=1;
   60084: out<=0;
   60085: out<=0;
   60086: out<=1;
   60087: out<=1;
   60088: out<=0;
   60089: out<=0;
   60090: out<=0;
   60091: out<=0;
   60092: out<=0;
   60093: out<=1;
   60094: out<=1;
   60095: out<=0;
   60096: out<=1;
   60097: out<=0;
   60098: out<=1;
   60099: out<=0;
   60100: out<=1;
   60101: out<=1;
   60102: out<=0;
   60103: out<=0;
   60104: out<=1;
   60105: out<=1;
   60106: out<=1;
   60107: out<=1;
   60108: out<=1;
   60109: out<=0;
   60110: out<=0;
   60111: out<=1;
   60112: out<=0;
   60113: out<=1;
   60114: out<=0;
   60115: out<=1;
   60116: out<=0;
   60117: out<=0;
   60118: out<=1;
   60119: out<=1;
   60120: out<=0;
   60121: out<=0;
   60122: out<=0;
   60123: out<=0;
   60124: out<=0;
   60125: out<=1;
   60126: out<=1;
   60127: out<=0;
   60128: out<=1;
   60129: out<=0;
   60130: out<=1;
   60131: out<=0;
   60132: out<=1;
   60133: out<=1;
   60134: out<=0;
   60135: out<=0;
   60136: out<=1;
   60137: out<=1;
   60138: out<=1;
   60139: out<=1;
   60140: out<=1;
   60141: out<=0;
   60142: out<=0;
   60143: out<=1;
   60144: out<=0;
   60145: out<=1;
   60146: out<=0;
   60147: out<=1;
   60148: out<=0;
   60149: out<=0;
   60150: out<=1;
   60151: out<=1;
   60152: out<=0;
   60153: out<=0;
   60154: out<=0;
   60155: out<=0;
   60156: out<=0;
   60157: out<=1;
   60158: out<=1;
   60159: out<=0;
   60160: out<=0;
   60161: out<=0;
   60162: out<=1;
   60163: out<=1;
   60164: out<=1;
   60165: out<=0;
   60166: out<=1;
   60167: out<=0;
   60168: out<=1;
   60169: out<=0;
   60170: out<=0;
   60171: out<=1;
   60172: out<=0;
   60173: out<=0;
   60174: out<=0;
   60175: out<=0;
   60176: out<=0;
   60177: out<=0;
   60178: out<=1;
   60179: out<=1;
   60180: out<=1;
   60181: out<=0;
   60182: out<=1;
   60183: out<=0;
   60184: out<=1;
   60185: out<=0;
   60186: out<=0;
   60187: out<=1;
   60188: out<=0;
   60189: out<=0;
   60190: out<=0;
   60191: out<=0;
   60192: out<=0;
   60193: out<=0;
   60194: out<=1;
   60195: out<=1;
   60196: out<=1;
   60197: out<=0;
   60198: out<=1;
   60199: out<=0;
   60200: out<=1;
   60201: out<=0;
   60202: out<=0;
   60203: out<=1;
   60204: out<=0;
   60205: out<=0;
   60206: out<=0;
   60207: out<=0;
   60208: out<=0;
   60209: out<=0;
   60210: out<=1;
   60211: out<=1;
   60212: out<=1;
   60213: out<=0;
   60214: out<=1;
   60215: out<=0;
   60216: out<=1;
   60217: out<=0;
   60218: out<=0;
   60219: out<=1;
   60220: out<=0;
   60221: out<=0;
   60222: out<=0;
   60223: out<=0;
   60224: out<=0;
   60225: out<=0;
   60226: out<=1;
   60227: out<=1;
   60228: out<=1;
   60229: out<=0;
   60230: out<=1;
   60231: out<=0;
   60232: out<=1;
   60233: out<=0;
   60234: out<=0;
   60235: out<=1;
   60236: out<=0;
   60237: out<=0;
   60238: out<=0;
   60239: out<=0;
   60240: out<=1;
   60241: out<=1;
   60242: out<=0;
   60243: out<=0;
   60244: out<=0;
   60245: out<=1;
   60246: out<=0;
   60247: out<=1;
   60248: out<=0;
   60249: out<=1;
   60250: out<=1;
   60251: out<=0;
   60252: out<=1;
   60253: out<=1;
   60254: out<=1;
   60255: out<=1;
   60256: out<=1;
   60257: out<=1;
   60258: out<=0;
   60259: out<=0;
   60260: out<=0;
   60261: out<=1;
   60262: out<=0;
   60263: out<=1;
   60264: out<=0;
   60265: out<=1;
   60266: out<=1;
   60267: out<=0;
   60268: out<=1;
   60269: out<=1;
   60270: out<=1;
   60271: out<=1;
   60272: out<=0;
   60273: out<=0;
   60274: out<=1;
   60275: out<=1;
   60276: out<=1;
   60277: out<=0;
   60278: out<=1;
   60279: out<=0;
   60280: out<=1;
   60281: out<=0;
   60282: out<=0;
   60283: out<=1;
   60284: out<=0;
   60285: out<=0;
   60286: out<=0;
   60287: out<=0;
   60288: out<=0;
   60289: out<=0;
   60290: out<=1;
   60291: out<=1;
   60292: out<=1;
   60293: out<=0;
   60294: out<=1;
   60295: out<=0;
   60296: out<=1;
   60297: out<=0;
   60298: out<=0;
   60299: out<=1;
   60300: out<=0;
   60301: out<=0;
   60302: out<=0;
   60303: out<=0;
   60304: out<=1;
   60305: out<=1;
   60306: out<=0;
   60307: out<=0;
   60308: out<=0;
   60309: out<=1;
   60310: out<=0;
   60311: out<=1;
   60312: out<=0;
   60313: out<=1;
   60314: out<=1;
   60315: out<=0;
   60316: out<=1;
   60317: out<=1;
   60318: out<=1;
   60319: out<=1;
   60320: out<=0;
   60321: out<=0;
   60322: out<=1;
   60323: out<=1;
   60324: out<=1;
   60325: out<=0;
   60326: out<=1;
   60327: out<=0;
   60328: out<=1;
   60329: out<=0;
   60330: out<=0;
   60331: out<=1;
   60332: out<=0;
   60333: out<=0;
   60334: out<=0;
   60335: out<=0;
   60336: out<=1;
   60337: out<=1;
   60338: out<=0;
   60339: out<=0;
   60340: out<=0;
   60341: out<=1;
   60342: out<=0;
   60343: out<=1;
   60344: out<=0;
   60345: out<=1;
   60346: out<=1;
   60347: out<=0;
   60348: out<=1;
   60349: out<=1;
   60350: out<=1;
   60351: out<=1;
   60352: out<=0;
   60353: out<=0;
   60354: out<=1;
   60355: out<=1;
   60356: out<=1;
   60357: out<=0;
   60358: out<=1;
   60359: out<=0;
   60360: out<=1;
   60361: out<=0;
   60362: out<=0;
   60363: out<=1;
   60364: out<=0;
   60365: out<=0;
   60366: out<=0;
   60367: out<=0;
   60368: out<=0;
   60369: out<=0;
   60370: out<=1;
   60371: out<=1;
   60372: out<=1;
   60373: out<=0;
   60374: out<=1;
   60375: out<=0;
   60376: out<=1;
   60377: out<=0;
   60378: out<=0;
   60379: out<=1;
   60380: out<=0;
   60381: out<=0;
   60382: out<=0;
   60383: out<=0;
   60384: out<=1;
   60385: out<=1;
   60386: out<=0;
   60387: out<=0;
   60388: out<=0;
   60389: out<=1;
   60390: out<=0;
   60391: out<=1;
   60392: out<=0;
   60393: out<=1;
   60394: out<=1;
   60395: out<=0;
   60396: out<=1;
   60397: out<=1;
   60398: out<=1;
   60399: out<=1;
   60400: out<=1;
   60401: out<=1;
   60402: out<=0;
   60403: out<=0;
   60404: out<=0;
   60405: out<=1;
   60406: out<=0;
   60407: out<=1;
   60408: out<=0;
   60409: out<=1;
   60410: out<=1;
   60411: out<=0;
   60412: out<=1;
   60413: out<=1;
   60414: out<=1;
   60415: out<=1;
   60416: out<=1;
   60417: out<=0;
   60418: out<=0;
   60419: out<=1;
   60420: out<=0;
   60421: out<=0;
   60422: out<=0;
   60423: out<=0;
   60424: out<=1;
   60425: out<=1;
   60426: out<=0;
   60427: out<=0;
   60428: out<=0;
   60429: out<=1;
   60430: out<=0;
   60431: out<=1;
   60432: out<=1;
   60433: out<=0;
   60434: out<=0;
   60435: out<=1;
   60436: out<=0;
   60437: out<=0;
   60438: out<=0;
   60439: out<=0;
   60440: out<=1;
   60441: out<=1;
   60442: out<=0;
   60443: out<=0;
   60444: out<=0;
   60445: out<=1;
   60446: out<=0;
   60447: out<=1;
   60448: out<=0;
   60449: out<=1;
   60450: out<=1;
   60451: out<=0;
   60452: out<=1;
   60453: out<=1;
   60454: out<=1;
   60455: out<=1;
   60456: out<=0;
   60457: out<=0;
   60458: out<=1;
   60459: out<=1;
   60460: out<=1;
   60461: out<=0;
   60462: out<=1;
   60463: out<=0;
   60464: out<=0;
   60465: out<=1;
   60466: out<=1;
   60467: out<=0;
   60468: out<=1;
   60469: out<=1;
   60470: out<=1;
   60471: out<=1;
   60472: out<=0;
   60473: out<=0;
   60474: out<=1;
   60475: out<=1;
   60476: out<=1;
   60477: out<=0;
   60478: out<=1;
   60479: out<=0;
   60480: out<=1;
   60481: out<=0;
   60482: out<=0;
   60483: out<=1;
   60484: out<=0;
   60485: out<=0;
   60486: out<=0;
   60487: out<=0;
   60488: out<=1;
   60489: out<=1;
   60490: out<=0;
   60491: out<=0;
   60492: out<=0;
   60493: out<=1;
   60494: out<=0;
   60495: out<=1;
   60496: out<=0;
   60497: out<=1;
   60498: out<=1;
   60499: out<=0;
   60500: out<=1;
   60501: out<=1;
   60502: out<=1;
   60503: out<=1;
   60504: out<=0;
   60505: out<=0;
   60506: out<=1;
   60507: out<=1;
   60508: out<=1;
   60509: out<=0;
   60510: out<=1;
   60511: out<=0;
   60512: out<=1;
   60513: out<=0;
   60514: out<=0;
   60515: out<=1;
   60516: out<=0;
   60517: out<=0;
   60518: out<=0;
   60519: out<=0;
   60520: out<=1;
   60521: out<=1;
   60522: out<=0;
   60523: out<=0;
   60524: out<=0;
   60525: out<=1;
   60526: out<=0;
   60527: out<=1;
   60528: out<=0;
   60529: out<=1;
   60530: out<=1;
   60531: out<=0;
   60532: out<=1;
   60533: out<=1;
   60534: out<=1;
   60535: out<=1;
   60536: out<=0;
   60537: out<=0;
   60538: out<=1;
   60539: out<=1;
   60540: out<=1;
   60541: out<=0;
   60542: out<=1;
   60543: out<=0;
   60544: out<=1;
   60545: out<=0;
   60546: out<=0;
   60547: out<=1;
   60548: out<=0;
   60549: out<=0;
   60550: out<=0;
   60551: out<=0;
   60552: out<=1;
   60553: out<=1;
   60554: out<=0;
   60555: out<=0;
   60556: out<=0;
   60557: out<=1;
   60558: out<=0;
   60559: out<=1;
   60560: out<=0;
   60561: out<=1;
   60562: out<=1;
   60563: out<=0;
   60564: out<=1;
   60565: out<=1;
   60566: out<=1;
   60567: out<=1;
   60568: out<=0;
   60569: out<=0;
   60570: out<=1;
   60571: out<=1;
   60572: out<=1;
   60573: out<=0;
   60574: out<=1;
   60575: out<=0;
   60576: out<=0;
   60577: out<=1;
   60578: out<=1;
   60579: out<=0;
   60580: out<=1;
   60581: out<=1;
   60582: out<=1;
   60583: out<=1;
   60584: out<=0;
   60585: out<=0;
   60586: out<=1;
   60587: out<=1;
   60588: out<=1;
   60589: out<=0;
   60590: out<=1;
   60591: out<=0;
   60592: out<=1;
   60593: out<=0;
   60594: out<=0;
   60595: out<=1;
   60596: out<=0;
   60597: out<=0;
   60598: out<=0;
   60599: out<=0;
   60600: out<=1;
   60601: out<=1;
   60602: out<=0;
   60603: out<=0;
   60604: out<=0;
   60605: out<=1;
   60606: out<=0;
   60607: out<=1;
   60608: out<=1;
   60609: out<=0;
   60610: out<=0;
   60611: out<=1;
   60612: out<=0;
   60613: out<=0;
   60614: out<=0;
   60615: out<=0;
   60616: out<=1;
   60617: out<=1;
   60618: out<=0;
   60619: out<=0;
   60620: out<=0;
   60621: out<=1;
   60622: out<=0;
   60623: out<=1;
   60624: out<=1;
   60625: out<=0;
   60626: out<=0;
   60627: out<=1;
   60628: out<=0;
   60629: out<=0;
   60630: out<=0;
   60631: out<=0;
   60632: out<=1;
   60633: out<=1;
   60634: out<=0;
   60635: out<=0;
   60636: out<=0;
   60637: out<=1;
   60638: out<=0;
   60639: out<=1;
   60640: out<=1;
   60641: out<=0;
   60642: out<=0;
   60643: out<=1;
   60644: out<=0;
   60645: out<=0;
   60646: out<=0;
   60647: out<=0;
   60648: out<=1;
   60649: out<=1;
   60650: out<=0;
   60651: out<=0;
   60652: out<=0;
   60653: out<=1;
   60654: out<=0;
   60655: out<=1;
   60656: out<=1;
   60657: out<=0;
   60658: out<=0;
   60659: out<=1;
   60660: out<=0;
   60661: out<=0;
   60662: out<=0;
   60663: out<=0;
   60664: out<=1;
   60665: out<=1;
   60666: out<=0;
   60667: out<=0;
   60668: out<=0;
   60669: out<=1;
   60670: out<=0;
   60671: out<=1;
   60672: out<=1;
   60673: out<=1;
   60674: out<=1;
   60675: out<=1;
   60676: out<=1;
   60677: out<=0;
   60678: out<=0;
   60679: out<=1;
   60680: out<=0;
   60681: out<=1;
   60682: out<=0;
   60683: out<=1;
   60684: out<=0;
   60685: out<=0;
   60686: out<=1;
   60687: out<=1;
   60688: out<=0;
   60689: out<=0;
   60690: out<=0;
   60691: out<=0;
   60692: out<=0;
   60693: out<=1;
   60694: out<=1;
   60695: out<=0;
   60696: out<=1;
   60697: out<=0;
   60698: out<=1;
   60699: out<=0;
   60700: out<=1;
   60701: out<=1;
   60702: out<=0;
   60703: out<=0;
   60704: out<=1;
   60705: out<=1;
   60706: out<=1;
   60707: out<=1;
   60708: out<=1;
   60709: out<=0;
   60710: out<=0;
   60711: out<=1;
   60712: out<=0;
   60713: out<=1;
   60714: out<=0;
   60715: out<=1;
   60716: out<=0;
   60717: out<=0;
   60718: out<=1;
   60719: out<=1;
   60720: out<=0;
   60721: out<=0;
   60722: out<=0;
   60723: out<=0;
   60724: out<=0;
   60725: out<=1;
   60726: out<=1;
   60727: out<=0;
   60728: out<=1;
   60729: out<=0;
   60730: out<=1;
   60731: out<=0;
   60732: out<=1;
   60733: out<=1;
   60734: out<=0;
   60735: out<=0;
   60736: out<=1;
   60737: out<=1;
   60738: out<=1;
   60739: out<=1;
   60740: out<=1;
   60741: out<=0;
   60742: out<=0;
   60743: out<=1;
   60744: out<=0;
   60745: out<=1;
   60746: out<=0;
   60747: out<=1;
   60748: out<=0;
   60749: out<=0;
   60750: out<=1;
   60751: out<=1;
   60752: out<=1;
   60753: out<=1;
   60754: out<=1;
   60755: out<=1;
   60756: out<=1;
   60757: out<=0;
   60758: out<=0;
   60759: out<=1;
   60760: out<=0;
   60761: out<=1;
   60762: out<=0;
   60763: out<=1;
   60764: out<=0;
   60765: out<=0;
   60766: out<=1;
   60767: out<=1;
   60768: out<=0;
   60769: out<=0;
   60770: out<=0;
   60771: out<=0;
   60772: out<=0;
   60773: out<=1;
   60774: out<=1;
   60775: out<=0;
   60776: out<=1;
   60777: out<=0;
   60778: out<=1;
   60779: out<=0;
   60780: out<=1;
   60781: out<=1;
   60782: out<=0;
   60783: out<=0;
   60784: out<=0;
   60785: out<=0;
   60786: out<=0;
   60787: out<=0;
   60788: out<=0;
   60789: out<=1;
   60790: out<=1;
   60791: out<=0;
   60792: out<=1;
   60793: out<=0;
   60794: out<=1;
   60795: out<=0;
   60796: out<=1;
   60797: out<=1;
   60798: out<=0;
   60799: out<=0;
   60800: out<=1;
   60801: out<=1;
   60802: out<=1;
   60803: out<=1;
   60804: out<=1;
   60805: out<=0;
   60806: out<=0;
   60807: out<=1;
   60808: out<=0;
   60809: out<=1;
   60810: out<=0;
   60811: out<=1;
   60812: out<=0;
   60813: out<=0;
   60814: out<=1;
   60815: out<=1;
   60816: out<=1;
   60817: out<=1;
   60818: out<=1;
   60819: out<=1;
   60820: out<=1;
   60821: out<=0;
   60822: out<=0;
   60823: out<=1;
   60824: out<=0;
   60825: out<=1;
   60826: out<=0;
   60827: out<=1;
   60828: out<=0;
   60829: out<=0;
   60830: out<=1;
   60831: out<=1;
   60832: out<=1;
   60833: out<=1;
   60834: out<=1;
   60835: out<=1;
   60836: out<=1;
   60837: out<=0;
   60838: out<=0;
   60839: out<=1;
   60840: out<=0;
   60841: out<=1;
   60842: out<=0;
   60843: out<=1;
   60844: out<=0;
   60845: out<=0;
   60846: out<=1;
   60847: out<=1;
   60848: out<=1;
   60849: out<=1;
   60850: out<=1;
   60851: out<=1;
   60852: out<=1;
   60853: out<=0;
   60854: out<=0;
   60855: out<=1;
   60856: out<=0;
   60857: out<=1;
   60858: out<=0;
   60859: out<=1;
   60860: out<=0;
   60861: out<=0;
   60862: out<=1;
   60863: out<=1;
   60864: out<=1;
   60865: out<=1;
   60866: out<=1;
   60867: out<=1;
   60868: out<=1;
   60869: out<=0;
   60870: out<=0;
   60871: out<=1;
   60872: out<=0;
   60873: out<=1;
   60874: out<=0;
   60875: out<=1;
   60876: out<=0;
   60877: out<=0;
   60878: out<=1;
   60879: out<=1;
   60880: out<=0;
   60881: out<=0;
   60882: out<=0;
   60883: out<=0;
   60884: out<=0;
   60885: out<=1;
   60886: out<=1;
   60887: out<=0;
   60888: out<=1;
   60889: out<=0;
   60890: out<=1;
   60891: out<=0;
   60892: out<=1;
   60893: out<=1;
   60894: out<=0;
   60895: out<=0;
   60896: out<=0;
   60897: out<=0;
   60898: out<=0;
   60899: out<=0;
   60900: out<=0;
   60901: out<=1;
   60902: out<=1;
   60903: out<=0;
   60904: out<=1;
   60905: out<=0;
   60906: out<=1;
   60907: out<=0;
   60908: out<=1;
   60909: out<=1;
   60910: out<=0;
   60911: out<=0;
   60912: out<=1;
   60913: out<=1;
   60914: out<=1;
   60915: out<=1;
   60916: out<=1;
   60917: out<=0;
   60918: out<=0;
   60919: out<=1;
   60920: out<=0;
   60921: out<=1;
   60922: out<=0;
   60923: out<=1;
   60924: out<=0;
   60925: out<=0;
   60926: out<=1;
   60927: out<=1;
   60928: out<=0;
   60929: out<=0;
   60930: out<=1;
   60931: out<=1;
   60932: out<=0;
   60933: out<=1;
   60934: out<=0;
   60935: out<=1;
   60936: out<=0;
   60937: out<=1;
   60938: out<=1;
   60939: out<=0;
   60940: out<=0;
   60941: out<=0;
   60942: out<=0;
   60943: out<=0;
   60944: out<=1;
   60945: out<=1;
   60946: out<=0;
   60947: out<=0;
   60948: out<=1;
   60949: out<=0;
   60950: out<=1;
   60951: out<=0;
   60952: out<=1;
   60953: out<=0;
   60954: out<=0;
   60955: out<=1;
   60956: out<=1;
   60957: out<=1;
   60958: out<=1;
   60959: out<=1;
   60960: out<=1;
   60961: out<=1;
   60962: out<=0;
   60963: out<=0;
   60964: out<=1;
   60965: out<=0;
   60966: out<=1;
   60967: out<=0;
   60968: out<=1;
   60969: out<=0;
   60970: out<=0;
   60971: out<=1;
   60972: out<=1;
   60973: out<=1;
   60974: out<=1;
   60975: out<=1;
   60976: out<=0;
   60977: out<=0;
   60978: out<=1;
   60979: out<=1;
   60980: out<=0;
   60981: out<=1;
   60982: out<=0;
   60983: out<=1;
   60984: out<=0;
   60985: out<=1;
   60986: out<=1;
   60987: out<=0;
   60988: out<=0;
   60989: out<=0;
   60990: out<=0;
   60991: out<=0;
   60992: out<=0;
   60993: out<=0;
   60994: out<=1;
   60995: out<=1;
   60996: out<=0;
   60997: out<=1;
   60998: out<=0;
   60999: out<=1;
   61000: out<=0;
   61001: out<=1;
   61002: out<=1;
   61003: out<=0;
   61004: out<=0;
   61005: out<=0;
   61006: out<=0;
   61007: out<=0;
   61008: out<=0;
   61009: out<=0;
   61010: out<=1;
   61011: out<=1;
   61012: out<=0;
   61013: out<=1;
   61014: out<=0;
   61015: out<=1;
   61016: out<=0;
   61017: out<=1;
   61018: out<=1;
   61019: out<=0;
   61020: out<=0;
   61021: out<=0;
   61022: out<=0;
   61023: out<=0;
   61024: out<=0;
   61025: out<=0;
   61026: out<=1;
   61027: out<=1;
   61028: out<=0;
   61029: out<=1;
   61030: out<=0;
   61031: out<=1;
   61032: out<=0;
   61033: out<=1;
   61034: out<=1;
   61035: out<=0;
   61036: out<=0;
   61037: out<=0;
   61038: out<=0;
   61039: out<=0;
   61040: out<=0;
   61041: out<=0;
   61042: out<=1;
   61043: out<=1;
   61044: out<=0;
   61045: out<=1;
   61046: out<=0;
   61047: out<=1;
   61048: out<=0;
   61049: out<=1;
   61050: out<=1;
   61051: out<=0;
   61052: out<=0;
   61053: out<=0;
   61054: out<=0;
   61055: out<=0;
   61056: out<=0;
   61057: out<=0;
   61058: out<=1;
   61059: out<=1;
   61060: out<=0;
   61061: out<=1;
   61062: out<=0;
   61063: out<=1;
   61064: out<=0;
   61065: out<=1;
   61066: out<=1;
   61067: out<=0;
   61068: out<=0;
   61069: out<=0;
   61070: out<=0;
   61071: out<=0;
   61072: out<=0;
   61073: out<=0;
   61074: out<=1;
   61075: out<=1;
   61076: out<=0;
   61077: out<=1;
   61078: out<=0;
   61079: out<=1;
   61080: out<=0;
   61081: out<=1;
   61082: out<=1;
   61083: out<=0;
   61084: out<=0;
   61085: out<=0;
   61086: out<=0;
   61087: out<=0;
   61088: out<=1;
   61089: out<=1;
   61090: out<=0;
   61091: out<=0;
   61092: out<=1;
   61093: out<=0;
   61094: out<=1;
   61095: out<=0;
   61096: out<=1;
   61097: out<=0;
   61098: out<=0;
   61099: out<=1;
   61100: out<=1;
   61101: out<=1;
   61102: out<=1;
   61103: out<=1;
   61104: out<=1;
   61105: out<=1;
   61106: out<=0;
   61107: out<=0;
   61108: out<=1;
   61109: out<=0;
   61110: out<=1;
   61111: out<=0;
   61112: out<=1;
   61113: out<=0;
   61114: out<=0;
   61115: out<=1;
   61116: out<=1;
   61117: out<=1;
   61118: out<=1;
   61119: out<=1;
   61120: out<=0;
   61121: out<=0;
   61122: out<=1;
   61123: out<=1;
   61124: out<=0;
   61125: out<=1;
   61126: out<=0;
   61127: out<=1;
   61128: out<=0;
   61129: out<=1;
   61130: out<=1;
   61131: out<=0;
   61132: out<=0;
   61133: out<=0;
   61134: out<=0;
   61135: out<=0;
   61136: out<=1;
   61137: out<=1;
   61138: out<=0;
   61139: out<=0;
   61140: out<=1;
   61141: out<=0;
   61142: out<=1;
   61143: out<=0;
   61144: out<=1;
   61145: out<=0;
   61146: out<=0;
   61147: out<=1;
   61148: out<=1;
   61149: out<=1;
   61150: out<=1;
   61151: out<=1;
   61152: out<=0;
   61153: out<=0;
   61154: out<=1;
   61155: out<=1;
   61156: out<=0;
   61157: out<=1;
   61158: out<=0;
   61159: out<=1;
   61160: out<=0;
   61161: out<=1;
   61162: out<=1;
   61163: out<=0;
   61164: out<=0;
   61165: out<=0;
   61166: out<=0;
   61167: out<=0;
   61168: out<=1;
   61169: out<=1;
   61170: out<=0;
   61171: out<=0;
   61172: out<=1;
   61173: out<=0;
   61174: out<=1;
   61175: out<=0;
   61176: out<=1;
   61177: out<=0;
   61178: out<=0;
   61179: out<=1;
   61180: out<=1;
   61181: out<=1;
   61182: out<=1;
   61183: out<=1;
   61184: out<=0;
   61185: out<=1;
   61186: out<=0;
   61187: out<=1;
   61188: out<=1;
   61189: out<=1;
   61190: out<=0;
   61191: out<=0;
   61192: out<=1;
   61193: out<=1;
   61194: out<=1;
   61195: out<=1;
   61196: out<=0;
   61197: out<=1;
   61198: out<=1;
   61199: out<=0;
   61200: out<=0;
   61201: out<=1;
   61202: out<=0;
   61203: out<=1;
   61204: out<=1;
   61205: out<=1;
   61206: out<=0;
   61207: out<=0;
   61208: out<=1;
   61209: out<=1;
   61210: out<=1;
   61211: out<=1;
   61212: out<=0;
   61213: out<=1;
   61214: out<=1;
   61215: out<=0;
   61216: out<=0;
   61217: out<=1;
   61218: out<=0;
   61219: out<=1;
   61220: out<=1;
   61221: out<=1;
   61222: out<=0;
   61223: out<=0;
   61224: out<=1;
   61225: out<=1;
   61226: out<=1;
   61227: out<=1;
   61228: out<=0;
   61229: out<=1;
   61230: out<=1;
   61231: out<=0;
   61232: out<=0;
   61233: out<=1;
   61234: out<=0;
   61235: out<=1;
   61236: out<=1;
   61237: out<=1;
   61238: out<=0;
   61239: out<=0;
   61240: out<=1;
   61241: out<=1;
   61242: out<=1;
   61243: out<=1;
   61244: out<=0;
   61245: out<=1;
   61246: out<=1;
   61247: out<=0;
   61248: out<=0;
   61249: out<=1;
   61250: out<=0;
   61251: out<=1;
   61252: out<=1;
   61253: out<=1;
   61254: out<=0;
   61255: out<=0;
   61256: out<=1;
   61257: out<=1;
   61258: out<=1;
   61259: out<=1;
   61260: out<=0;
   61261: out<=1;
   61262: out<=1;
   61263: out<=0;
   61264: out<=1;
   61265: out<=0;
   61266: out<=1;
   61267: out<=0;
   61268: out<=0;
   61269: out<=0;
   61270: out<=1;
   61271: out<=1;
   61272: out<=0;
   61273: out<=0;
   61274: out<=0;
   61275: out<=0;
   61276: out<=1;
   61277: out<=0;
   61278: out<=0;
   61279: out<=1;
   61280: out<=1;
   61281: out<=0;
   61282: out<=1;
   61283: out<=0;
   61284: out<=0;
   61285: out<=0;
   61286: out<=1;
   61287: out<=1;
   61288: out<=0;
   61289: out<=0;
   61290: out<=0;
   61291: out<=0;
   61292: out<=1;
   61293: out<=0;
   61294: out<=0;
   61295: out<=1;
   61296: out<=0;
   61297: out<=1;
   61298: out<=0;
   61299: out<=1;
   61300: out<=1;
   61301: out<=1;
   61302: out<=0;
   61303: out<=0;
   61304: out<=1;
   61305: out<=1;
   61306: out<=1;
   61307: out<=1;
   61308: out<=0;
   61309: out<=1;
   61310: out<=1;
   61311: out<=0;
   61312: out<=0;
   61313: out<=1;
   61314: out<=0;
   61315: out<=1;
   61316: out<=1;
   61317: out<=1;
   61318: out<=0;
   61319: out<=0;
   61320: out<=1;
   61321: out<=1;
   61322: out<=1;
   61323: out<=1;
   61324: out<=0;
   61325: out<=1;
   61326: out<=1;
   61327: out<=0;
   61328: out<=1;
   61329: out<=0;
   61330: out<=1;
   61331: out<=0;
   61332: out<=0;
   61333: out<=0;
   61334: out<=1;
   61335: out<=1;
   61336: out<=0;
   61337: out<=0;
   61338: out<=0;
   61339: out<=0;
   61340: out<=1;
   61341: out<=0;
   61342: out<=0;
   61343: out<=1;
   61344: out<=0;
   61345: out<=1;
   61346: out<=0;
   61347: out<=1;
   61348: out<=1;
   61349: out<=1;
   61350: out<=0;
   61351: out<=0;
   61352: out<=1;
   61353: out<=1;
   61354: out<=1;
   61355: out<=1;
   61356: out<=0;
   61357: out<=1;
   61358: out<=1;
   61359: out<=0;
   61360: out<=1;
   61361: out<=0;
   61362: out<=1;
   61363: out<=0;
   61364: out<=0;
   61365: out<=0;
   61366: out<=1;
   61367: out<=1;
   61368: out<=0;
   61369: out<=0;
   61370: out<=0;
   61371: out<=0;
   61372: out<=1;
   61373: out<=0;
   61374: out<=0;
   61375: out<=1;
   61376: out<=0;
   61377: out<=1;
   61378: out<=0;
   61379: out<=1;
   61380: out<=1;
   61381: out<=1;
   61382: out<=0;
   61383: out<=0;
   61384: out<=1;
   61385: out<=1;
   61386: out<=1;
   61387: out<=1;
   61388: out<=0;
   61389: out<=1;
   61390: out<=1;
   61391: out<=0;
   61392: out<=0;
   61393: out<=1;
   61394: out<=0;
   61395: out<=1;
   61396: out<=1;
   61397: out<=1;
   61398: out<=0;
   61399: out<=0;
   61400: out<=1;
   61401: out<=1;
   61402: out<=1;
   61403: out<=1;
   61404: out<=0;
   61405: out<=1;
   61406: out<=1;
   61407: out<=0;
   61408: out<=1;
   61409: out<=0;
   61410: out<=1;
   61411: out<=0;
   61412: out<=0;
   61413: out<=0;
   61414: out<=1;
   61415: out<=1;
   61416: out<=0;
   61417: out<=0;
   61418: out<=0;
   61419: out<=0;
   61420: out<=1;
   61421: out<=0;
   61422: out<=0;
   61423: out<=1;
   61424: out<=1;
   61425: out<=0;
   61426: out<=1;
   61427: out<=0;
   61428: out<=0;
   61429: out<=0;
   61430: out<=1;
   61431: out<=1;
   61432: out<=0;
   61433: out<=0;
   61434: out<=0;
   61435: out<=0;
   61436: out<=1;
   61437: out<=0;
   61438: out<=0;
   61439: out<=1;
   61440: out<=1;
   61441: out<=1;
   61442: out<=0;
   61443: out<=0;
   61444: out<=0;
   61445: out<=1;
   61446: out<=0;
   61447: out<=1;
   61448: out<=1;
   61449: out<=0;
   61450: out<=0;
   61451: out<=1;
   61452: out<=0;
   61453: out<=0;
   61454: out<=0;
   61455: out<=0;
   61456: out<=0;
   61457: out<=0;
   61458: out<=1;
   61459: out<=1;
   61460: out<=1;
   61461: out<=0;
   61462: out<=1;
   61463: out<=0;
   61464: out<=0;
   61465: out<=1;
   61466: out<=1;
   61467: out<=0;
   61468: out<=1;
   61469: out<=1;
   61470: out<=1;
   61471: out<=1;
   61472: out<=1;
   61473: out<=1;
   61474: out<=0;
   61475: out<=0;
   61476: out<=0;
   61477: out<=1;
   61478: out<=0;
   61479: out<=1;
   61480: out<=1;
   61481: out<=0;
   61482: out<=0;
   61483: out<=1;
   61484: out<=0;
   61485: out<=0;
   61486: out<=0;
   61487: out<=0;
   61488: out<=0;
   61489: out<=0;
   61490: out<=1;
   61491: out<=1;
   61492: out<=1;
   61493: out<=0;
   61494: out<=1;
   61495: out<=0;
   61496: out<=0;
   61497: out<=1;
   61498: out<=1;
   61499: out<=0;
   61500: out<=1;
   61501: out<=1;
   61502: out<=1;
   61503: out<=1;
   61504: out<=0;
   61505: out<=0;
   61506: out<=1;
   61507: out<=1;
   61508: out<=1;
   61509: out<=0;
   61510: out<=1;
   61511: out<=0;
   61512: out<=0;
   61513: out<=1;
   61514: out<=1;
   61515: out<=0;
   61516: out<=1;
   61517: out<=1;
   61518: out<=1;
   61519: out<=1;
   61520: out<=0;
   61521: out<=0;
   61522: out<=1;
   61523: out<=1;
   61524: out<=1;
   61525: out<=0;
   61526: out<=1;
   61527: out<=0;
   61528: out<=0;
   61529: out<=1;
   61530: out<=1;
   61531: out<=0;
   61532: out<=1;
   61533: out<=1;
   61534: out<=1;
   61535: out<=1;
   61536: out<=1;
   61537: out<=1;
   61538: out<=0;
   61539: out<=0;
   61540: out<=0;
   61541: out<=1;
   61542: out<=0;
   61543: out<=1;
   61544: out<=1;
   61545: out<=0;
   61546: out<=0;
   61547: out<=1;
   61548: out<=0;
   61549: out<=0;
   61550: out<=0;
   61551: out<=0;
   61552: out<=1;
   61553: out<=1;
   61554: out<=0;
   61555: out<=0;
   61556: out<=0;
   61557: out<=1;
   61558: out<=0;
   61559: out<=1;
   61560: out<=1;
   61561: out<=0;
   61562: out<=0;
   61563: out<=1;
   61564: out<=0;
   61565: out<=0;
   61566: out<=0;
   61567: out<=0;
   61568: out<=0;
   61569: out<=0;
   61570: out<=1;
   61571: out<=1;
   61572: out<=1;
   61573: out<=0;
   61574: out<=1;
   61575: out<=0;
   61576: out<=0;
   61577: out<=1;
   61578: out<=1;
   61579: out<=0;
   61580: out<=1;
   61581: out<=1;
   61582: out<=1;
   61583: out<=1;
   61584: out<=0;
   61585: out<=0;
   61586: out<=1;
   61587: out<=1;
   61588: out<=1;
   61589: out<=0;
   61590: out<=1;
   61591: out<=0;
   61592: out<=0;
   61593: out<=1;
   61594: out<=1;
   61595: out<=0;
   61596: out<=1;
   61597: out<=1;
   61598: out<=1;
   61599: out<=1;
   61600: out<=0;
   61601: out<=0;
   61602: out<=1;
   61603: out<=1;
   61604: out<=1;
   61605: out<=0;
   61606: out<=1;
   61607: out<=0;
   61608: out<=0;
   61609: out<=1;
   61610: out<=1;
   61611: out<=0;
   61612: out<=1;
   61613: out<=1;
   61614: out<=1;
   61615: out<=1;
   61616: out<=0;
   61617: out<=0;
   61618: out<=1;
   61619: out<=1;
   61620: out<=1;
   61621: out<=0;
   61622: out<=1;
   61623: out<=0;
   61624: out<=0;
   61625: out<=1;
   61626: out<=1;
   61627: out<=0;
   61628: out<=1;
   61629: out<=1;
   61630: out<=1;
   61631: out<=1;
   61632: out<=1;
   61633: out<=1;
   61634: out<=0;
   61635: out<=0;
   61636: out<=0;
   61637: out<=1;
   61638: out<=0;
   61639: out<=1;
   61640: out<=1;
   61641: out<=0;
   61642: out<=0;
   61643: out<=1;
   61644: out<=0;
   61645: out<=0;
   61646: out<=0;
   61647: out<=0;
   61648: out<=0;
   61649: out<=0;
   61650: out<=1;
   61651: out<=1;
   61652: out<=1;
   61653: out<=0;
   61654: out<=1;
   61655: out<=0;
   61656: out<=0;
   61657: out<=1;
   61658: out<=1;
   61659: out<=0;
   61660: out<=1;
   61661: out<=1;
   61662: out<=1;
   61663: out<=1;
   61664: out<=0;
   61665: out<=0;
   61666: out<=1;
   61667: out<=1;
   61668: out<=1;
   61669: out<=0;
   61670: out<=1;
   61671: out<=0;
   61672: out<=0;
   61673: out<=1;
   61674: out<=1;
   61675: out<=0;
   61676: out<=1;
   61677: out<=1;
   61678: out<=1;
   61679: out<=1;
   61680: out<=1;
   61681: out<=1;
   61682: out<=0;
   61683: out<=0;
   61684: out<=0;
   61685: out<=1;
   61686: out<=0;
   61687: out<=1;
   61688: out<=1;
   61689: out<=0;
   61690: out<=0;
   61691: out<=1;
   61692: out<=0;
   61693: out<=0;
   61694: out<=0;
   61695: out<=0;
   61696: out<=1;
   61697: out<=0;
   61698: out<=1;
   61699: out<=0;
   61700: out<=1;
   61701: out<=1;
   61702: out<=0;
   61703: out<=0;
   61704: out<=0;
   61705: out<=0;
   61706: out<=0;
   61707: out<=0;
   61708: out<=0;
   61709: out<=1;
   61710: out<=1;
   61711: out<=0;
   61712: out<=1;
   61713: out<=0;
   61714: out<=1;
   61715: out<=0;
   61716: out<=1;
   61717: out<=1;
   61718: out<=0;
   61719: out<=0;
   61720: out<=0;
   61721: out<=0;
   61722: out<=0;
   61723: out<=0;
   61724: out<=0;
   61725: out<=1;
   61726: out<=1;
   61727: out<=0;
   61728: out<=0;
   61729: out<=1;
   61730: out<=0;
   61731: out<=1;
   61732: out<=0;
   61733: out<=0;
   61734: out<=1;
   61735: out<=1;
   61736: out<=1;
   61737: out<=1;
   61738: out<=1;
   61739: out<=1;
   61740: out<=1;
   61741: out<=0;
   61742: out<=0;
   61743: out<=1;
   61744: out<=0;
   61745: out<=1;
   61746: out<=0;
   61747: out<=1;
   61748: out<=0;
   61749: out<=0;
   61750: out<=1;
   61751: out<=1;
   61752: out<=1;
   61753: out<=1;
   61754: out<=1;
   61755: out<=1;
   61756: out<=1;
   61757: out<=0;
   61758: out<=0;
   61759: out<=1;
   61760: out<=0;
   61761: out<=1;
   61762: out<=0;
   61763: out<=1;
   61764: out<=0;
   61765: out<=0;
   61766: out<=1;
   61767: out<=1;
   61768: out<=1;
   61769: out<=1;
   61770: out<=1;
   61771: out<=1;
   61772: out<=1;
   61773: out<=0;
   61774: out<=0;
   61775: out<=1;
   61776: out<=1;
   61777: out<=0;
   61778: out<=1;
   61779: out<=0;
   61780: out<=1;
   61781: out<=1;
   61782: out<=0;
   61783: out<=0;
   61784: out<=0;
   61785: out<=0;
   61786: out<=0;
   61787: out<=0;
   61788: out<=0;
   61789: out<=1;
   61790: out<=1;
   61791: out<=0;
   61792: out<=0;
   61793: out<=1;
   61794: out<=0;
   61795: out<=1;
   61796: out<=0;
   61797: out<=0;
   61798: out<=1;
   61799: out<=1;
   61800: out<=1;
   61801: out<=1;
   61802: out<=1;
   61803: out<=1;
   61804: out<=1;
   61805: out<=0;
   61806: out<=0;
   61807: out<=1;
   61808: out<=1;
   61809: out<=0;
   61810: out<=1;
   61811: out<=0;
   61812: out<=1;
   61813: out<=1;
   61814: out<=0;
   61815: out<=0;
   61816: out<=0;
   61817: out<=0;
   61818: out<=0;
   61819: out<=0;
   61820: out<=0;
   61821: out<=1;
   61822: out<=1;
   61823: out<=0;
   61824: out<=0;
   61825: out<=1;
   61826: out<=0;
   61827: out<=1;
   61828: out<=0;
   61829: out<=0;
   61830: out<=1;
   61831: out<=1;
   61832: out<=1;
   61833: out<=1;
   61834: out<=1;
   61835: out<=1;
   61836: out<=1;
   61837: out<=0;
   61838: out<=0;
   61839: out<=1;
   61840: out<=1;
   61841: out<=0;
   61842: out<=1;
   61843: out<=0;
   61844: out<=1;
   61845: out<=1;
   61846: out<=0;
   61847: out<=0;
   61848: out<=0;
   61849: out<=0;
   61850: out<=0;
   61851: out<=0;
   61852: out<=0;
   61853: out<=1;
   61854: out<=1;
   61855: out<=0;
   61856: out<=1;
   61857: out<=0;
   61858: out<=1;
   61859: out<=0;
   61860: out<=1;
   61861: out<=1;
   61862: out<=0;
   61863: out<=0;
   61864: out<=0;
   61865: out<=0;
   61866: out<=0;
   61867: out<=0;
   61868: out<=0;
   61869: out<=1;
   61870: out<=1;
   61871: out<=0;
   61872: out<=0;
   61873: out<=1;
   61874: out<=0;
   61875: out<=1;
   61876: out<=0;
   61877: out<=0;
   61878: out<=1;
   61879: out<=1;
   61880: out<=1;
   61881: out<=1;
   61882: out<=1;
   61883: out<=1;
   61884: out<=1;
   61885: out<=0;
   61886: out<=0;
   61887: out<=1;
   61888: out<=1;
   61889: out<=0;
   61890: out<=1;
   61891: out<=0;
   61892: out<=1;
   61893: out<=1;
   61894: out<=0;
   61895: out<=0;
   61896: out<=0;
   61897: out<=0;
   61898: out<=0;
   61899: out<=0;
   61900: out<=0;
   61901: out<=1;
   61902: out<=1;
   61903: out<=0;
   61904: out<=1;
   61905: out<=0;
   61906: out<=1;
   61907: out<=0;
   61908: out<=1;
   61909: out<=1;
   61910: out<=0;
   61911: out<=0;
   61912: out<=0;
   61913: out<=0;
   61914: out<=0;
   61915: out<=0;
   61916: out<=0;
   61917: out<=1;
   61918: out<=1;
   61919: out<=0;
   61920: out<=1;
   61921: out<=0;
   61922: out<=1;
   61923: out<=0;
   61924: out<=1;
   61925: out<=1;
   61926: out<=0;
   61927: out<=0;
   61928: out<=0;
   61929: out<=0;
   61930: out<=0;
   61931: out<=0;
   61932: out<=0;
   61933: out<=1;
   61934: out<=1;
   61935: out<=0;
   61936: out<=1;
   61937: out<=0;
   61938: out<=1;
   61939: out<=0;
   61940: out<=1;
   61941: out<=1;
   61942: out<=0;
   61943: out<=0;
   61944: out<=0;
   61945: out<=0;
   61946: out<=0;
   61947: out<=0;
   61948: out<=0;
   61949: out<=1;
   61950: out<=1;
   61951: out<=0;
   61952: out<=1;
   61953: out<=0;
   61954: out<=0;
   61955: out<=1;
   61956: out<=1;
   61957: out<=1;
   61958: out<=1;
   61959: out<=1;
   61960: out<=1;
   61961: out<=1;
   61962: out<=0;
   61963: out<=0;
   61964: out<=1;
   61965: out<=0;
   61966: out<=1;
   61967: out<=0;
   61968: out<=1;
   61969: out<=0;
   61970: out<=0;
   61971: out<=1;
   61972: out<=1;
   61973: out<=1;
   61974: out<=1;
   61975: out<=1;
   61976: out<=1;
   61977: out<=1;
   61978: out<=0;
   61979: out<=0;
   61980: out<=1;
   61981: out<=0;
   61982: out<=1;
   61983: out<=0;
   61984: out<=1;
   61985: out<=0;
   61986: out<=0;
   61987: out<=1;
   61988: out<=1;
   61989: out<=1;
   61990: out<=1;
   61991: out<=1;
   61992: out<=1;
   61993: out<=1;
   61994: out<=0;
   61995: out<=0;
   61996: out<=1;
   61997: out<=0;
   61998: out<=1;
   61999: out<=0;
   62000: out<=1;
   62001: out<=0;
   62002: out<=0;
   62003: out<=1;
   62004: out<=1;
   62005: out<=1;
   62006: out<=1;
   62007: out<=1;
   62008: out<=1;
   62009: out<=1;
   62010: out<=0;
   62011: out<=0;
   62012: out<=1;
   62013: out<=0;
   62014: out<=1;
   62015: out<=0;
   62016: out<=0;
   62017: out<=1;
   62018: out<=1;
   62019: out<=0;
   62020: out<=0;
   62021: out<=0;
   62022: out<=0;
   62023: out<=0;
   62024: out<=0;
   62025: out<=0;
   62026: out<=1;
   62027: out<=1;
   62028: out<=0;
   62029: out<=1;
   62030: out<=0;
   62031: out<=1;
   62032: out<=1;
   62033: out<=0;
   62034: out<=0;
   62035: out<=1;
   62036: out<=1;
   62037: out<=1;
   62038: out<=1;
   62039: out<=1;
   62040: out<=1;
   62041: out<=1;
   62042: out<=0;
   62043: out<=0;
   62044: out<=1;
   62045: out<=0;
   62046: out<=1;
   62047: out<=0;
   62048: out<=1;
   62049: out<=0;
   62050: out<=0;
   62051: out<=1;
   62052: out<=1;
   62053: out<=1;
   62054: out<=1;
   62055: out<=1;
   62056: out<=1;
   62057: out<=1;
   62058: out<=0;
   62059: out<=0;
   62060: out<=1;
   62061: out<=0;
   62062: out<=1;
   62063: out<=0;
   62064: out<=0;
   62065: out<=1;
   62066: out<=1;
   62067: out<=0;
   62068: out<=0;
   62069: out<=0;
   62070: out<=0;
   62071: out<=0;
   62072: out<=0;
   62073: out<=0;
   62074: out<=1;
   62075: out<=1;
   62076: out<=0;
   62077: out<=1;
   62078: out<=0;
   62079: out<=1;
   62080: out<=0;
   62081: out<=1;
   62082: out<=1;
   62083: out<=0;
   62084: out<=0;
   62085: out<=0;
   62086: out<=0;
   62087: out<=0;
   62088: out<=0;
   62089: out<=0;
   62090: out<=1;
   62091: out<=1;
   62092: out<=0;
   62093: out<=1;
   62094: out<=0;
   62095: out<=1;
   62096: out<=1;
   62097: out<=0;
   62098: out<=0;
   62099: out<=1;
   62100: out<=1;
   62101: out<=1;
   62102: out<=1;
   62103: out<=1;
   62104: out<=1;
   62105: out<=1;
   62106: out<=0;
   62107: out<=0;
   62108: out<=1;
   62109: out<=0;
   62110: out<=1;
   62111: out<=0;
   62112: out<=0;
   62113: out<=1;
   62114: out<=1;
   62115: out<=0;
   62116: out<=0;
   62117: out<=0;
   62118: out<=0;
   62119: out<=0;
   62120: out<=0;
   62121: out<=0;
   62122: out<=1;
   62123: out<=1;
   62124: out<=0;
   62125: out<=1;
   62126: out<=0;
   62127: out<=1;
   62128: out<=1;
   62129: out<=0;
   62130: out<=0;
   62131: out<=1;
   62132: out<=1;
   62133: out<=1;
   62134: out<=1;
   62135: out<=1;
   62136: out<=1;
   62137: out<=1;
   62138: out<=0;
   62139: out<=0;
   62140: out<=1;
   62141: out<=0;
   62142: out<=1;
   62143: out<=0;
   62144: out<=1;
   62145: out<=0;
   62146: out<=0;
   62147: out<=1;
   62148: out<=1;
   62149: out<=1;
   62150: out<=1;
   62151: out<=1;
   62152: out<=1;
   62153: out<=1;
   62154: out<=0;
   62155: out<=0;
   62156: out<=1;
   62157: out<=0;
   62158: out<=1;
   62159: out<=0;
   62160: out<=1;
   62161: out<=0;
   62162: out<=0;
   62163: out<=1;
   62164: out<=1;
   62165: out<=1;
   62166: out<=1;
   62167: out<=1;
   62168: out<=1;
   62169: out<=1;
   62170: out<=0;
   62171: out<=0;
   62172: out<=1;
   62173: out<=0;
   62174: out<=1;
   62175: out<=0;
   62176: out<=0;
   62177: out<=1;
   62178: out<=1;
   62179: out<=0;
   62180: out<=0;
   62181: out<=0;
   62182: out<=0;
   62183: out<=0;
   62184: out<=0;
   62185: out<=0;
   62186: out<=1;
   62187: out<=1;
   62188: out<=0;
   62189: out<=1;
   62190: out<=0;
   62191: out<=1;
   62192: out<=0;
   62193: out<=1;
   62194: out<=1;
   62195: out<=0;
   62196: out<=0;
   62197: out<=0;
   62198: out<=0;
   62199: out<=0;
   62200: out<=0;
   62201: out<=0;
   62202: out<=1;
   62203: out<=1;
   62204: out<=0;
   62205: out<=1;
   62206: out<=0;
   62207: out<=1;
   62208: out<=1;
   62209: out<=1;
   62210: out<=1;
   62211: out<=1;
   62212: out<=0;
   62213: out<=1;
   62214: out<=1;
   62215: out<=0;
   62216: out<=0;
   62217: out<=1;
   62218: out<=0;
   62219: out<=1;
   62220: out<=1;
   62221: out<=1;
   62222: out<=0;
   62223: out<=0;
   62224: out<=0;
   62225: out<=0;
   62226: out<=0;
   62227: out<=0;
   62228: out<=1;
   62229: out<=0;
   62230: out<=0;
   62231: out<=1;
   62232: out<=1;
   62233: out<=0;
   62234: out<=1;
   62235: out<=0;
   62236: out<=0;
   62237: out<=0;
   62238: out<=1;
   62239: out<=1;
   62240: out<=0;
   62241: out<=0;
   62242: out<=0;
   62243: out<=0;
   62244: out<=1;
   62245: out<=0;
   62246: out<=0;
   62247: out<=1;
   62248: out<=1;
   62249: out<=0;
   62250: out<=1;
   62251: out<=0;
   62252: out<=0;
   62253: out<=0;
   62254: out<=1;
   62255: out<=1;
   62256: out<=1;
   62257: out<=1;
   62258: out<=1;
   62259: out<=1;
   62260: out<=0;
   62261: out<=1;
   62262: out<=1;
   62263: out<=0;
   62264: out<=0;
   62265: out<=1;
   62266: out<=0;
   62267: out<=1;
   62268: out<=1;
   62269: out<=1;
   62270: out<=0;
   62271: out<=0;
   62272: out<=0;
   62273: out<=0;
   62274: out<=0;
   62275: out<=0;
   62276: out<=1;
   62277: out<=0;
   62278: out<=0;
   62279: out<=1;
   62280: out<=1;
   62281: out<=0;
   62282: out<=1;
   62283: out<=0;
   62284: out<=0;
   62285: out<=0;
   62286: out<=1;
   62287: out<=1;
   62288: out<=0;
   62289: out<=0;
   62290: out<=0;
   62291: out<=0;
   62292: out<=1;
   62293: out<=0;
   62294: out<=0;
   62295: out<=1;
   62296: out<=1;
   62297: out<=0;
   62298: out<=1;
   62299: out<=0;
   62300: out<=0;
   62301: out<=0;
   62302: out<=1;
   62303: out<=1;
   62304: out<=0;
   62305: out<=0;
   62306: out<=0;
   62307: out<=0;
   62308: out<=1;
   62309: out<=0;
   62310: out<=0;
   62311: out<=1;
   62312: out<=1;
   62313: out<=0;
   62314: out<=1;
   62315: out<=0;
   62316: out<=0;
   62317: out<=0;
   62318: out<=1;
   62319: out<=1;
   62320: out<=0;
   62321: out<=0;
   62322: out<=0;
   62323: out<=0;
   62324: out<=1;
   62325: out<=0;
   62326: out<=0;
   62327: out<=1;
   62328: out<=1;
   62329: out<=0;
   62330: out<=1;
   62331: out<=0;
   62332: out<=0;
   62333: out<=0;
   62334: out<=1;
   62335: out<=1;
   62336: out<=0;
   62337: out<=0;
   62338: out<=0;
   62339: out<=0;
   62340: out<=1;
   62341: out<=0;
   62342: out<=0;
   62343: out<=1;
   62344: out<=1;
   62345: out<=0;
   62346: out<=1;
   62347: out<=0;
   62348: out<=0;
   62349: out<=0;
   62350: out<=1;
   62351: out<=1;
   62352: out<=0;
   62353: out<=0;
   62354: out<=0;
   62355: out<=0;
   62356: out<=1;
   62357: out<=0;
   62358: out<=0;
   62359: out<=1;
   62360: out<=1;
   62361: out<=0;
   62362: out<=1;
   62363: out<=0;
   62364: out<=0;
   62365: out<=0;
   62366: out<=1;
   62367: out<=1;
   62368: out<=1;
   62369: out<=1;
   62370: out<=1;
   62371: out<=1;
   62372: out<=0;
   62373: out<=1;
   62374: out<=1;
   62375: out<=0;
   62376: out<=0;
   62377: out<=1;
   62378: out<=0;
   62379: out<=1;
   62380: out<=1;
   62381: out<=1;
   62382: out<=0;
   62383: out<=0;
   62384: out<=1;
   62385: out<=1;
   62386: out<=1;
   62387: out<=1;
   62388: out<=0;
   62389: out<=1;
   62390: out<=1;
   62391: out<=0;
   62392: out<=0;
   62393: out<=1;
   62394: out<=0;
   62395: out<=1;
   62396: out<=1;
   62397: out<=1;
   62398: out<=0;
   62399: out<=0;
   62400: out<=1;
   62401: out<=1;
   62402: out<=1;
   62403: out<=1;
   62404: out<=0;
   62405: out<=1;
   62406: out<=1;
   62407: out<=0;
   62408: out<=0;
   62409: out<=1;
   62410: out<=0;
   62411: out<=1;
   62412: out<=1;
   62413: out<=1;
   62414: out<=0;
   62415: out<=0;
   62416: out<=0;
   62417: out<=0;
   62418: out<=0;
   62419: out<=0;
   62420: out<=1;
   62421: out<=0;
   62422: out<=0;
   62423: out<=1;
   62424: out<=1;
   62425: out<=0;
   62426: out<=1;
   62427: out<=0;
   62428: out<=0;
   62429: out<=0;
   62430: out<=1;
   62431: out<=1;
   62432: out<=1;
   62433: out<=1;
   62434: out<=1;
   62435: out<=1;
   62436: out<=0;
   62437: out<=1;
   62438: out<=1;
   62439: out<=0;
   62440: out<=0;
   62441: out<=1;
   62442: out<=0;
   62443: out<=1;
   62444: out<=1;
   62445: out<=1;
   62446: out<=0;
   62447: out<=0;
   62448: out<=0;
   62449: out<=0;
   62450: out<=0;
   62451: out<=0;
   62452: out<=1;
   62453: out<=0;
   62454: out<=0;
   62455: out<=1;
   62456: out<=1;
   62457: out<=0;
   62458: out<=1;
   62459: out<=0;
   62460: out<=0;
   62461: out<=0;
   62462: out<=1;
   62463: out<=1;
   62464: out<=1;
   62465: out<=0;
   62466: out<=1;
   62467: out<=0;
   62468: out<=0;
   62469: out<=0;
   62470: out<=1;
   62471: out<=1;
   62472: out<=1;
   62473: out<=1;
   62474: out<=1;
   62475: out<=1;
   62476: out<=0;
   62477: out<=1;
   62478: out<=1;
   62479: out<=0;
   62480: out<=0;
   62481: out<=1;
   62482: out<=0;
   62483: out<=1;
   62484: out<=1;
   62485: out<=1;
   62486: out<=0;
   62487: out<=0;
   62488: out<=0;
   62489: out<=0;
   62490: out<=0;
   62491: out<=0;
   62492: out<=1;
   62493: out<=0;
   62494: out<=0;
   62495: out<=1;
   62496: out<=1;
   62497: out<=0;
   62498: out<=1;
   62499: out<=0;
   62500: out<=0;
   62501: out<=0;
   62502: out<=1;
   62503: out<=1;
   62504: out<=1;
   62505: out<=1;
   62506: out<=1;
   62507: out<=1;
   62508: out<=0;
   62509: out<=1;
   62510: out<=1;
   62511: out<=0;
   62512: out<=0;
   62513: out<=1;
   62514: out<=0;
   62515: out<=1;
   62516: out<=1;
   62517: out<=1;
   62518: out<=0;
   62519: out<=0;
   62520: out<=0;
   62521: out<=0;
   62522: out<=0;
   62523: out<=0;
   62524: out<=1;
   62525: out<=0;
   62526: out<=0;
   62527: out<=1;
   62528: out<=0;
   62529: out<=1;
   62530: out<=0;
   62531: out<=1;
   62532: out<=1;
   62533: out<=1;
   62534: out<=0;
   62535: out<=0;
   62536: out<=0;
   62537: out<=0;
   62538: out<=0;
   62539: out<=0;
   62540: out<=1;
   62541: out<=0;
   62542: out<=0;
   62543: out<=1;
   62544: out<=0;
   62545: out<=1;
   62546: out<=0;
   62547: out<=1;
   62548: out<=1;
   62549: out<=1;
   62550: out<=0;
   62551: out<=0;
   62552: out<=0;
   62553: out<=0;
   62554: out<=0;
   62555: out<=0;
   62556: out<=1;
   62557: out<=0;
   62558: out<=0;
   62559: out<=1;
   62560: out<=1;
   62561: out<=0;
   62562: out<=1;
   62563: out<=0;
   62564: out<=0;
   62565: out<=0;
   62566: out<=1;
   62567: out<=1;
   62568: out<=1;
   62569: out<=1;
   62570: out<=1;
   62571: out<=1;
   62572: out<=0;
   62573: out<=1;
   62574: out<=1;
   62575: out<=0;
   62576: out<=1;
   62577: out<=0;
   62578: out<=1;
   62579: out<=0;
   62580: out<=0;
   62581: out<=0;
   62582: out<=1;
   62583: out<=1;
   62584: out<=1;
   62585: out<=1;
   62586: out<=1;
   62587: out<=1;
   62588: out<=0;
   62589: out<=1;
   62590: out<=1;
   62591: out<=0;
   62592: out<=0;
   62593: out<=1;
   62594: out<=0;
   62595: out<=1;
   62596: out<=1;
   62597: out<=1;
   62598: out<=0;
   62599: out<=0;
   62600: out<=0;
   62601: out<=0;
   62602: out<=0;
   62603: out<=0;
   62604: out<=1;
   62605: out<=0;
   62606: out<=0;
   62607: out<=1;
   62608: out<=0;
   62609: out<=1;
   62610: out<=0;
   62611: out<=1;
   62612: out<=1;
   62613: out<=1;
   62614: out<=0;
   62615: out<=0;
   62616: out<=0;
   62617: out<=0;
   62618: out<=0;
   62619: out<=0;
   62620: out<=1;
   62621: out<=0;
   62622: out<=0;
   62623: out<=1;
   62624: out<=0;
   62625: out<=1;
   62626: out<=0;
   62627: out<=1;
   62628: out<=1;
   62629: out<=1;
   62630: out<=0;
   62631: out<=0;
   62632: out<=0;
   62633: out<=0;
   62634: out<=0;
   62635: out<=0;
   62636: out<=1;
   62637: out<=0;
   62638: out<=0;
   62639: out<=1;
   62640: out<=0;
   62641: out<=1;
   62642: out<=0;
   62643: out<=1;
   62644: out<=1;
   62645: out<=1;
   62646: out<=0;
   62647: out<=0;
   62648: out<=0;
   62649: out<=0;
   62650: out<=0;
   62651: out<=0;
   62652: out<=1;
   62653: out<=0;
   62654: out<=0;
   62655: out<=1;
   62656: out<=1;
   62657: out<=0;
   62658: out<=1;
   62659: out<=0;
   62660: out<=0;
   62661: out<=0;
   62662: out<=1;
   62663: out<=1;
   62664: out<=1;
   62665: out<=1;
   62666: out<=1;
   62667: out<=1;
   62668: out<=0;
   62669: out<=1;
   62670: out<=1;
   62671: out<=0;
   62672: out<=0;
   62673: out<=1;
   62674: out<=0;
   62675: out<=1;
   62676: out<=1;
   62677: out<=1;
   62678: out<=0;
   62679: out<=0;
   62680: out<=0;
   62681: out<=0;
   62682: out<=0;
   62683: out<=0;
   62684: out<=1;
   62685: out<=0;
   62686: out<=0;
   62687: out<=1;
   62688: out<=0;
   62689: out<=1;
   62690: out<=0;
   62691: out<=1;
   62692: out<=1;
   62693: out<=1;
   62694: out<=0;
   62695: out<=0;
   62696: out<=0;
   62697: out<=0;
   62698: out<=0;
   62699: out<=0;
   62700: out<=1;
   62701: out<=0;
   62702: out<=0;
   62703: out<=1;
   62704: out<=1;
   62705: out<=0;
   62706: out<=1;
   62707: out<=0;
   62708: out<=0;
   62709: out<=0;
   62710: out<=1;
   62711: out<=1;
   62712: out<=1;
   62713: out<=1;
   62714: out<=1;
   62715: out<=1;
   62716: out<=0;
   62717: out<=1;
   62718: out<=1;
   62719: out<=0;
   62720: out<=0;
   62721: out<=0;
   62722: out<=1;
   62723: out<=1;
   62724: out<=0;
   62725: out<=1;
   62726: out<=0;
   62727: out<=1;
   62728: out<=1;
   62729: out<=0;
   62730: out<=0;
   62731: out<=1;
   62732: out<=1;
   62733: out<=1;
   62734: out<=1;
   62735: out<=1;
   62736: out<=0;
   62737: out<=0;
   62738: out<=1;
   62739: out<=1;
   62740: out<=0;
   62741: out<=1;
   62742: out<=0;
   62743: out<=1;
   62744: out<=1;
   62745: out<=0;
   62746: out<=0;
   62747: out<=1;
   62748: out<=1;
   62749: out<=1;
   62750: out<=1;
   62751: out<=1;
   62752: out<=1;
   62753: out<=1;
   62754: out<=0;
   62755: out<=0;
   62756: out<=1;
   62757: out<=0;
   62758: out<=1;
   62759: out<=0;
   62760: out<=0;
   62761: out<=1;
   62762: out<=1;
   62763: out<=0;
   62764: out<=0;
   62765: out<=0;
   62766: out<=0;
   62767: out<=0;
   62768: out<=1;
   62769: out<=1;
   62770: out<=0;
   62771: out<=0;
   62772: out<=1;
   62773: out<=0;
   62774: out<=1;
   62775: out<=0;
   62776: out<=0;
   62777: out<=1;
   62778: out<=1;
   62779: out<=0;
   62780: out<=0;
   62781: out<=0;
   62782: out<=0;
   62783: out<=0;
   62784: out<=1;
   62785: out<=1;
   62786: out<=0;
   62787: out<=0;
   62788: out<=1;
   62789: out<=0;
   62790: out<=1;
   62791: out<=0;
   62792: out<=0;
   62793: out<=1;
   62794: out<=1;
   62795: out<=0;
   62796: out<=0;
   62797: out<=0;
   62798: out<=0;
   62799: out<=0;
   62800: out<=0;
   62801: out<=0;
   62802: out<=1;
   62803: out<=1;
   62804: out<=0;
   62805: out<=1;
   62806: out<=0;
   62807: out<=1;
   62808: out<=1;
   62809: out<=0;
   62810: out<=0;
   62811: out<=1;
   62812: out<=1;
   62813: out<=1;
   62814: out<=1;
   62815: out<=1;
   62816: out<=1;
   62817: out<=1;
   62818: out<=0;
   62819: out<=0;
   62820: out<=1;
   62821: out<=0;
   62822: out<=1;
   62823: out<=0;
   62824: out<=0;
   62825: out<=1;
   62826: out<=1;
   62827: out<=0;
   62828: out<=0;
   62829: out<=0;
   62830: out<=0;
   62831: out<=0;
   62832: out<=0;
   62833: out<=0;
   62834: out<=1;
   62835: out<=1;
   62836: out<=0;
   62837: out<=1;
   62838: out<=0;
   62839: out<=1;
   62840: out<=1;
   62841: out<=0;
   62842: out<=0;
   62843: out<=1;
   62844: out<=1;
   62845: out<=1;
   62846: out<=1;
   62847: out<=1;
   62848: out<=1;
   62849: out<=1;
   62850: out<=0;
   62851: out<=0;
   62852: out<=1;
   62853: out<=0;
   62854: out<=1;
   62855: out<=0;
   62856: out<=0;
   62857: out<=1;
   62858: out<=1;
   62859: out<=0;
   62860: out<=0;
   62861: out<=0;
   62862: out<=0;
   62863: out<=0;
   62864: out<=0;
   62865: out<=0;
   62866: out<=1;
   62867: out<=1;
   62868: out<=0;
   62869: out<=1;
   62870: out<=0;
   62871: out<=1;
   62872: out<=1;
   62873: out<=0;
   62874: out<=0;
   62875: out<=1;
   62876: out<=1;
   62877: out<=1;
   62878: out<=1;
   62879: out<=1;
   62880: out<=0;
   62881: out<=0;
   62882: out<=1;
   62883: out<=1;
   62884: out<=0;
   62885: out<=1;
   62886: out<=0;
   62887: out<=1;
   62888: out<=1;
   62889: out<=0;
   62890: out<=0;
   62891: out<=1;
   62892: out<=1;
   62893: out<=1;
   62894: out<=1;
   62895: out<=1;
   62896: out<=1;
   62897: out<=1;
   62898: out<=0;
   62899: out<=0;
   62900: out<=1;
   62901: out<=0;
   62902: out<=1;
   62903: out<=0;
   62904: out<=0;
   62905: out<=1;
   62906: out<=1;
   62907: out<=0;
   62908: out<=0;
   62909: out<=0;
   62910: out<=0;
   62911: out<=0;
   62912: out<=0;
   62913: out<=0;
   62914: out<=1;
   62915: out<=1;
   62916: out<=0;
   62917: out<=1;
   62918: out<=0;
   62919: out<=1;
   62920: out<=1;
   62921: out<=0;
   62922: out<=0;
   62923: out<=1;
   62924: out<=1;
   62925: out<=1;
   62926: out<=1;
   62927: out<=1;
   62928: out<=0;
   62929: out<=0;
   62930: out<=1;
   62931: out<=1;
   62932: out<=0;
   62933: out<=1;
   62934: out<=0;
   62935: out<=1;
   62936: out<=1;
   62937: out<=0;
   62938: out<=0;
   62939: out<=1;
   62940: out<=1;
   62941: out<=1;
   62942: out<=1;
   62943: out<=1;
   62944: out<=0;
   62945: out<=0;
   62946: out<=1;
   62947: out<=1;
   62948: out<=0;
   62949: out<=1;
   62950: out<=0;
   62951: out<=1;
   62952: out<=1;
   62953: out<=0;
   62954: out<=0;
   62955: out<=1;
   62956: out<=1;
   62957: out<=1;
   62958: out<=1;
   62959: out<=1;
   62960: out<=0;
   62961: out<=0;
   62962: out<=1;
   62963: out<=1;
   62964: out<=0;
   62965: out<=1;
   62966: out<=0;
   62967: out<=1;
   62968: out<=1;
   62969: out<=0;
   62970: out<=0;
   62971: out<=1;
   62972: out<=1;
   62973: out<=1;
   62974: out<=1;
   62975: out<=1;
   62976: out<=0;
   62977: out<=0;
   62978: out<=0;
   62979: out<=0;
   62980: out<=0;
   62981: out<=1;
   62982: out<=1;
   62983: out<=0;
   62984: out<=0;
   62985: out<=1;
   62986: out<=0;
   62987: out<=1;
   62988: out<=0;
   62989: out<=0;
   62990: out<=1;
   62991: out<=1;
   62992: out<=0;
   62993: out<=0;
   62994: out<=0;
   62995: out<=0;
   62996: out<=0;
   62997: out<=1;
   62998: out<=1;
   62999: out<=0;
   63000: out<=0;
   63001: out<=1;
   63002: out<=0;
   63003: out<=1;
   63004: out<=0;
   63005: out<=0;
   63006: out<=1;
   63007: out<=1;
   63008: out<=0;
   63009: out<=0;
   63010: out<=0;
   63011: out<=0;
   63012: out<=0;
   63013: out<=1;
   63014: out<=1;
   63015: out<=0;
   63016: out<=0;
   63017: out<=1;
   63018: out<=0;
   63019: out<=1;
   63020: out<=0;
   63021: out<=0;
   63022: out<=1;
   63023: out<=1;
   63024: out<=0;
   63025: out<=0;
   63026: out<=0;
   63027: out<=0;
   63028: out<=0;
   63029: out<=1;
   63030: out<=1;
   63031: out<=0;
   63032: out<=0;
   63033: out<=1;
   63034: out<=0;
   63035: out<=1;
   63036: out<=0;
   63037: out<=0;
   63038: out<=1;
   63039: out<=1;
   63040: out<=1;
   63041: out<=1;
   63042: out<=1;
   63043: out<=1;
   63044: out<=1;
   63045: out<=0;
   63046: out<=0;
   63047: out<=1;
   63048: out<=1;
   63049: out<=0;
   63050: out<=1;
   63051: out<=0;
   63052: out<=1;
   63053: out<=1;
   63054: out<=0;
   63055: out<=0;
   63056: out<=0;
   63057: out<=0;
   63058: out<=0;
   63059: out<=0;
   63060: out<=0;
   63061: out<=1;
   63062: out<=1;
   63063: out<=0;
   63064: out<=0;
   63065: out<=1;
   63066: out<=0;
   63067: out<=1;
   63068: out<=0;
   63069: out<=0;
   63070: out<=1;
   63071: out<=1;
   63072: out<=0;
   63073: out<=0;
   63074: out<=0;
   63075: out<=0;
   63076: out<=0;
   63077: out<=1;
   63078: out<=1;
   63079: out<=0;
   63080: out<=0;
   63081: out<=1;
   63082: out<=0;
   63083: out<=1;
   63084: out<=0;
   63085: out<=0;
   63086: out<=1;
   63087: out<=1;
   63088: out<=1;
   63089: out<=1;
   63090: out<=1;
   63091: out<=1;
   63092: out<=1;
   63093: out<=0;
   63094: out<=0;
   63095: out<=1;
   63096: out<=1;
   63097: out<=0;
   63098: out<=1;
   63099: out<=0;
   63100: out<=1;
   63101: out<=1;
   63102: out<=0;
   63103: out<=0;
   63104: out<=1;
   63105: out<=1;
   63106: out<=1;
   63107: out<=1;
   63108: out<=1;
   63109: out<=0;
   63110: out<=0;
   63111: out<=1;
   63112: out<=1;
   63113: out<=0;
   63114: out<=1;
   63115: out<=0;
   63116: out<=1;
   63117: out<=1;
   63118: out<=0;
   63119: out<=0;
   63120: out<=0;
   63121: out<=0;
   63122: out<=0;
   63123: out<=0;
   63124: out<=0;
   63125: out<=1;
   63126: out<=1;
   63127: out<=0;
   63128: out<=0;
   63129: out<=1;
   63130: out<=0;
   63131: out<=1;
   63132: out<=0;
   63133: out<=0;
   63134: out<=1;
   63135: out<=1;
   63136: out<=1;
   63137: out<=1;
   63138: out<=1;
   63139: out<=1;
   63140: out<=1;
   63141: out<=0;
   63142: out<=0;
   63143: out<=1;
   63144: out<=1;
   63145: out<=0;
   63146: out<=1;
   63147: out<=0;
   63148: out<=1;
   63149: out<=1;
   63150: out<=0;
   63151: out<=0;
   63152: out<=0;
   63153: out<=0;
   63154: out<=0;
   63155: out<=0;
   63156: out<=0;
   63157: out<=1;
   63158: out<=1;
   63159: out<=0;
   63160: out<=0;
   63161: out<=1;
   63162: out<=0;
   63163: out<=1;
   63164: out<=0;
   63165: out<=0;
   63166: out<=1;
   63167: out<=1;
   63168: out<=0;
   63169: out<=0;
   63170: out<=0;
   63171: out<=0;
   63172: out<=0;
   63173: out<=1;
   63174: out<=1;
   63175: out<=0;
   63176: out<=0;
   63177: out<=1;
   63178: out<=0;
   63179: out<=1;
   63180: out<=0;
   63181: out<=0;
   63182: out<=1;
   63183: out<=1;
   63184: out<=0;
   63185: out<=0;
   63186: out<=0;
   63187: out<=0;
   63188: out<=0;
   63189: out<=1;
   63190: out<=1;
   63191: out<=0;
   63192: out<=0;
   63193: out<=1;
   63194: out<=0;
   63195: out<=1;
   63196: out<=0;
   63197: out<=0;
   63198: out<=1;
   63199: out<=1;
   63200: out<=1;
   63201: out<=1;
   63202: out<=1;
   63203: out<=1;
   63204: out<=1;
   63205: out<=0;
   63206: out<=0;
   63207: out<=1;
   63208: out<=1;
   63209: out<=0;
   63210: out<=1;
   63211: out<=0;
   63212: out<=1;
   63213: out<=1;
   63214: out<=0;
   63215: out<=0;
   63216: out<=1;
   63217: out<=1;
   63218: out<=1;
   63219: out<=1;
   63220: out<=1;
   63221: out<=0;
   63222: out<=0;
   63223: out<=1;
   63224: out<=1;
   63225: out<=0;
   63226: out<=1;
   63227: out<=0;
   63228: out<=1;
   63229: out<=1;
   63230: out<=0;
   63231: out<=0;
   63232: out<=1;
   63233: out<=0;
   63234: out<=0;
   63235: out<=1;
   63236: out<=0;
   63237: out<=0;
   63238: out<=0;
   63239: out<=0;
   63240: out<=0;
   63241: out<=0;
   63242: out<=1;
   63243: out<=1;
   63244: out<=1;
   63245: out<=0;
   63246: out<=1;
   63247: out<=0;
   63248: out<=0;
   63249: out<=1;
   63250: out<=1;
   63251: out<=0;
   63252: out<=1;
   63253: out<=1;
   63254: out<=1;
   63255: out<=1;
   63256: out<=1;
   63257: out<=1;
   63258: out<=0;
   63259: out<=0;
   63260: out<=0;
   63261: out<=1;
   63262: out<=0;
   63263: out<=1;
   63264: out<=0;
   63265: out<=1;
   63266: out<=1;
   63267: out<=0;
   63268: out<=1;
   63269: out<=1;
   63270: out<=1;
   63271: out<=1;
   63272: out<=1;
   63273: out<=1;
   63274: out<=0;
   63275: out<=0;
   63276: out<=0;
   63277: out<=1;
   63278: out<=0;
   63279: out<=1;
   63280: out<=1;
   63281: out<=0;
   63282: out<=0;
   63283: out<=1;
   63284: out<=0;
   63285: out<=0;
   63286: out<=0;
   63287: out<=0;
   63288: out<=0;
   63289: out<=0;
   63290: out<=1;
   63291: out<=1;
   63292: out<=1;
   63293: out<=0;
   63294: out<=1;
   63295: out<=0;
   63296: out<=0;
   63297: out<=1;
   63298: out<=1;
   63299: out<=0;
   63300: out<=1;
   63301: out<=1;
   63302: out<=1;
   63303: out<=1;
   63304: out<=1;
   63305: out<=1;
   63306: out<=0;
   63307: out<=0;
   63308: out<=0;
   63309: out<=1;
   63310: out<=0;
   63311: out<=1;
   63312: out<=0;
   63313: out<=1;
   63314: out<=1;
   63315: out<=0;
   63316: out<=1;
   63317: out<=1;
   63318: out<=1;
   63319: out<=1;
   63320: out<=1;
   63321: out<=1;
   63322: out<=0;
   63323: out<=0;
   63324: out<=0;
   63325: out<=1;
   63326: out<=0;
   63327: out<=1;
   63328: out<=0;
   63329: out<=1;
   63330: out<=1;
   63331: out<=0;
   63332: out<=1;
   63333: out<=1;
   63334: out<=1;
   63335: out<=1;
   63336: out<=1;
   63337: out<=1;
   63338: out<=0;
   63339: out<=0;
   63340: out<=0;
   63341: out<=1;
   63342: out<=0;
   63343: out<=1;
   63344: out<=0;
   63345: out<=1;
   63346: out<=1;
   63347: out<=0;
   63348: out<=1;
   63349: out<=1;
   63350: out<=1;
   63351: out<=1;
   63352: out<=1;
   63353: out<=1;
   63354: out<=0;
   63355: out<=0;
   63356: out<=0;
   63357: out<=1;
   63358: out<=0;
   63359: out<=1;
   63360: out<=0;
   63361: out<=1;
   63362: out<=1;
   63363: out<=0;
   63364: out<=1;
   63365: out<=1;
   63366: out<=1;
   63367: out<=1;
   63368: out<=1;
   63369: out<=1;
   63370: out<=0;
   63371: out<=0;
   63372: out<=0;
   63373: out<=1;
   63374: out<=0;
   63375: out<=1;
   63376: out<=0;
   63377: out<=1;
   63378: out<=1;
   63379: out<=0;
   63380: out<=1;
   63381: out<=1;
   63382: out<=1;
   63383: out<=1;
   63384: out<=1;
   63385: out<=1;
   63386: out<=0;
   63387: out<=0;
   63388: out<=0;
   63389: out<=1;
   63390: out<=0;
   63391: out<=1;
   63392: out<=1;
   63393: out<=0;
   63394: out<=0;
   63395: out<=1;
   63396: out<=0;
   63397: out<=0;
   63398: out<=0;
   63399: out<=0;
   63400: out<=0;
   63401: out<=0;
   63402: out<=1;
   63403: out<=1;
   63404: out<=1;
   63405: out<=0;
   63406: out<=1;
   63407: out<=0;
   63408: out<=1;
   63409: out<=0;
   63410: out<=0;
   63411: out<=1;
   63412: out<=0;
   63413: out<=0;
   63414: out<=0;
   63415: out<=0;
   63416: out<=0;
   63417: out<=0;
   63418: out<=1;
   63419: out<=1;
   63420: out<=1;
   63421: out<=0;
   63422: out<=1;
   63423: out<=0;
   63424: out<=1;
   63425: out<=0;
   63426: out<=0;
   63427: out<=1;
   63428: out<=0;
   63429: out<=0;
   63430: out<=0;
   63431: out<=0;
   63432: out<=0;
   63433: out<=0;
   63434: out<=1;
   63435: out<=1;
   63436: out<=1;
   63437: out<=0;
   63438: out<=1;
   63439: out<=0;
   63440: out<=0;
   63441: out<=1;
   63442: out<=1;
   63443: out<=0;
   63444: out<=1;
   63445: out<=1;
   63446: out<=1;
   63447: out<=1;
   63448: out<=1;
   63449: out<=1;
   63450: out<=0;
   63451: out<=0;
   63452: out<=0;
   63453: out<=1;
   63454: out<=0;
   63455: out<=1;
   63456: out<=1;
   63457: out<=0;
   63458: out<=0;
   63459: out<=1;
   63460: out<=0;
   63461: out<=0;
   63462: out<=0;
   63463: out<=0;
   63464: out<=0;
   63465: out<=0;
   63466: out<=1;
   63467: out<=1;
   63468: out<=1;
   63469: out<=0;
   63470: out<=1;
   63471: out<=0;
   63472: out<=0;
   63473: out<=1;
   63474: out<=1;
   63475: out<=0;
   63476: out<=1;
   63477: out<=1;
   63478: out<=1;
   63479: out<=1;
   63480: out<=1;
   63481: out<=1;
   63482: out<=0;
   63483: out<=0;
   63484: out<=0;
   63485: out<=1;
   63486: out<=0;
   63487: out<=1;
   63488: out<=1;
   63489: out<=0;
   63490: out<=0;
   63491: out<=1;
   63492: out<=0;
   63493: out<=0;
   63494: out<=0;
   63495: out<=0;
   63496: out<=1;
   63497: out<=1;
   63498: out<=0;
   63499: out<=0;
   63500: out<=0;
   63501: out<=1;
   63502: out<=0;
   63503: out<=1;
   63504: out<=0;
   63505: out<=1;
   63506: out<=1;
   63507: out<=0;
   63508: out<=1;
   63509: out<=1;
   63510: out<=1;
   63511: out<=1;
   63512: out<=0;
   63513: out<=0;
   63514: out<=1;
   63515: out<=1;
   63516: out<=1;
   63517: out<=0;
   63518: out<=1;
   63519: out<=0;
   63520: out<=1;
   63521: out<=0;
   63522: out<=0;
   63523: out<=1;
   63524: out<=0;
   63525: out<=0;
   63526: out<=0;
   63527: out<=0;
   63528: out<=1;
   63529: out<=1;
   63530: out<=0;
   63531: out<=0;
   63532: out<=0;
   63533: out<=1;
   63534: out<=0;
   63535: out<=1;
   63536: out<=0;
   63537: out<=1;
   63538: out<=1;
   63539: out<=0;
   63540: out<=1;
   63541: out<=1;
   63542: out<=1;
   63543: out<=1;
   63544: out<=0;
   63545: out<=0;
   63546: out<=1;
   63547: out<=1;
   63548: out<=1;
   63549: out<=0;
   63550: out<=1;
   63551: out<=0;
   63552: out<=0;
   63553: out<=1;
   63554: out<=1;
   63555: out<=0;
   63556: out<=1;
   63557: out<=1;
   63558: out<=1;
   63559: out<=1;
   63560: out<=0;
   63561: out<=0;
   63562: out<=1;
   63563: out<=1;
   63564: out<=1;
   63565: out<=0;
   63566: out<=1;
   63567: out<=0;
   63568: out<=0;
   63569: out<=1;
   63570: out<=1;
   63571: out<=0;
   63572: out<=1;
   63573: out<=1;
   63574: out<=1;
   63575: out<=1;
   63576: out<=0;
   63577: out<=0;
   63578: out<=1;
   63579: out<=1;
   63580: out<=1;
   63581: out<=0;
   63582: out<=1;
   63583: out<=0;
   63584: out<=1;
   63585: out<=0;
   63586: out<=0;
   63587: out<=1;
   63588: out<=0;
   63589: out<=0;
   63590: out<=0;
   63591: out<=0;
   63592: out<=1;
   63593: out<=1;
   63594: out<=0;
   63595: out<=0;
   63596: out<=0;
   63597: out<=1;
   63598: out<=0;
   63599: out<=1;
   63600: out<=1;
   63601: out<=0;
   63602: out<=0;
   63603: out<=1;
   63604: out<=0;
   63605: out<=0;
   63606: out<=0;
   63607: out<=0;
   63608: out<=1;
   63609: out<=1;
   63610: out<=0;
   63611: out<=0;
   63612: out<=0;
   63613: out<=1;
   63614: out<=0;
   63615: out<=1;
   63616: out<=0;
   63617: out<=1;
   63618: out<=1;
   63619: out<=0;
   63620: out<=1;
   63621: out<=1;
   63622: out<=1;
   63623: out<=1;
   63624: out<=0;
   63625: out<=0;
   63626: out<=1;
   63627: out<=1;
   63628: out<=1;
   63629: out<=0;
   63630: out<=1;
   63631: out<=0;
   63632: out<=0;
   63633: out<=1;
   63634: out<=1;
   63635: out<=0;
   63636: out<=1;
   63637: out<=1;
   63638: out<=1;
   63639: out<=1;
   63640: out<=0;
   63641: out<=0;
   63642: out<=1;
   63643: out<=1;
   63644: out<=1;
   63645: out<=0;
   63646: out<=1;
   63647: out<=0;
   63648: out<=0;
   63649: out<=1;
   63650: out<=1;
   63651: out<=0;
   63652: out<=1;
   63653: out<=1;
   63654: out<=1;
   63655: out<=1;
   63656: out<=0;
   63657: out<=0;
   63658: out<=1;
   63659: out<=1;
   63660: out<=1;
   63661: out<=0;
   63662: out<=1;
   63663: out<=0;
   63664: out<=0;
   63665: out<=1;
   63666: out<=1;
   63667: out<=0;
   63668: out<=1;
   63669: out<=1;
   63670: out<=1;
   63671: out<=1;
   63672: out<=0;
   63673: out<=0;
   63674: out<=1;
   63675: out<=1;
   63676: out<=1;
   63677: out<=0;
   63678: out<=1;
   63679: out<=0;
   63680: out<=1;
   63681: out<=0;
   63682: out<=0;
   63683: out<=1;
   63684: out<=0;
   63685: out<=0;
   63686: out<=0;
   63687: out<=0;
   63688: out<=1;
   63689: out<=1;
   63690: out<=0;
   63691: out<=0;
   63692: out<=0;
   63693: out<=1;
   63694: out<=0;
   63695: out<=1;
   63696: out<=0;
   63697: out<=1;
   63698: out<=1;
   63699: out<=0;
   63700: out<=1;
   63701: out<=1;
   63702: out<=1;
   63703: out<=1;
   63704: out<=0;
   63705: out<=0;
   63706: out<=1;
   63707: out<=1;
   63708: out<=1;
   63709: out<=0;
   63710: out<=1;
   63711: out<=0;
   63712: out<=0;
   63713: out<=1;
   63714: out<=1;
   63715: out<=0;
   63716: out<=1;
   63717: out<=1;
   63718: out<=1;
   63719: out<=1;
   63720: out<=0;
   63721: out<=0;
   63722: out<=1;
   63723: out<=1;
   63724: out<=1;
   63725: out<=0;
   63726: out<=1;
   63727: out<=0;
   63728: out<=1;
   63729: out<=0;
   63730: out<=0;
   63731: out<=1;
   63732: out<=0;
   63733: out<=0;
   63734: out<=0;
   63735: out<=0;
   63736: out<=1;
   63737: out<=1;
   63738: out<=0;
   63739: out<=0;
   63740: out<=0;
   63741: out<=1;
   63742: out<=0;
   63743: out<=1;
   63744: out<=0;
   63745: out<=0;
   63746: out<=0;
   63747: out<=0;
   63748: out<=0;
   63749: out<=1;
   63750: out<=1;
   63751: out<=0;
   63752: out<=1;
   63753: out<=0;
   63754: out<=1;
   63755: out<=0;
   63756: out<=1;
   63757: out<=1;
   63758: out<=0;
   63759: out<=0;
   63760: out<=0;
   63761: out<=0;
   63762: out<=0;
   63763: out<=0;
   63764: out<=0;
   63765: out<=1;
   63766: out<=1;
   63767: out<=0;
   63768: out<=1;
   63769: out<=0;
   63770: out<=1;
   63771: out<=0;
   63772: out<=1;
   63773: out<=1;
   63774: out<=0;
   63775: out<=0;
   63776: out<=1;
   63777: out<=1;
   63778: out<=1;
   63779: out<=1;
   63780: out<=1;
   63781: out<=0;
   63782: out<=0;
   63783: out<=1;
   63784: out<=0;
   63785: out<=1;
   63786: out<=0;
   63787: out<=1;
   63788: out<=0;
   63789: out<=0;
   63790: out<=1;
   63791: out<=1;
   63792: out<=1;
   63793: out<=1;
   63794: out<=1;
   63795: out<=1;
   63796: out<=1;
   63797: out<=0;
   63798: out<=0;
   63799: out<=1;
   63800: out<=0;
   63801: out<=1;
   63802: out<=0;
   63803: out<=1;
   63804: out<=0;
   63805: out<=0;
   63806: out<=1;
   63807: out<=1;
   63808: out<=1;
   63809: out<=1;
   63810: out<=1;
   63811: out<=1;
   63812: out<=1;
   63813: out<=0;
   63814: out<=0;
   63815: out<=1;
   63816: out<=0;
   63817: out<=1;
   63818: out<=0;
   63819: out<=1;
   63820: out<=0;
   63821: out<=0;
   63822: out<=1;
   63823: out<=1;
   63824: out<=0;
   63825: out<=0;
   63826: out<=0;
   63827: out<=0;
   63828: out<=0;
   63829: out<=1;
   63830: out<=1;
   63831: out<=0;
   63832: out<=1;
   63833: out<=0;
   63834: out<=1;
   63835: out<=0;
   63836: out<=1;
   63837: out<=1;
   63838: out<=0;
   63839: out<=0;
   63840: out<=1;
   63841: out<=1;
   63842: out<=1;
   63843: out<=1;
   63844: out<=1;
   63845: out<=0;
   63846: out<=0;
   63847: out<=1;
   63848: out<=0;
   63849: out<=1;
   63850: out<=0;
   63851: out<=1;
   63852: out<=0;
   63853: out<=0;
   63854: out<=1;
   63855: out<=1;
   63856: out<=0;
   63857: out<=0;
   63858: out<=0;
   63859: out<=0;
   63860: out<=0;
   63861: out<=1;
   63862: out<=1;
   63863: out<=0;
   63864: out<=1;
   63865: out<=0;
   63866: out<=1;
   63867: out<=0;
   63868: out<=1;
   63869: out<=1;
   63870: out<=0;
   63871: out<=0;
   63872: out<=1;
   63873: out<=1;
   63874: out<=1;
   63875: out<=1;
   63876: out<=1;
   63877: out<=0;
   63878: out<=0;
   63879: out<=1;
   63880: out<=0;
   63881: out<=1;
   63882: out<=0;
   63883: out<=1;
   63884: out<=0;
   63885: out<=0;
   63886: out<=1;
   63887: out<=1;
   63888: out<=0;
   63889: out<=0;
   63890: out<=0;
   63891: out<=0;
   63892: out<=0;
   63893: out<=1;
   63894: out<=1;
   63895: out<=0;
   63896: out<=1;
   63897: out<=0;
   63898: out<=1;
   63899: out<=0;
   63900: out<=1;
   63901: out<=1;
   63902: out<=0;
   63903: out<=0;
   63904: out<=0;
   63905: out<=0;
   63906: out<=0;
   63907: out<=0;
   63908: out<=0;
   63909: out<=1;
   63910: out<=1;
   63911: out<=0;
   63912: out<=1;
   63913: out<=0;
   63914: out<=1;
   63915: out<=0;
   63916: out<=1;
   63917: out<=1;
   63918: out<=0;
   63919: out<=0;
   63920: out<=1;
   63921: out<=1;
   63922: out<=1;
   63923: out<=1;
   63924: out<=1;
   63925: out<=0;
   63926: out<=0;
   63927: out<=1;
   63928: out<=0;
   63929: out<=1;
   63930: out<=0;
   63931: out<=1;
   63932: out<=0;
   63933: out<=0;
   63934: out<=1;
   63935: out<=1;
   63936: out<=0;
   63937: out<=0;
   63938: out<=0;
   63939: out<=0;
   63940: out<=0;
   63941: out<=1;
   63942: out<=1;
   63943: out<=0;
   63944: out<=1;
   63945: out<=0;
   63946: out<=1;
   63947: out<=0;
   63948: out<=1;
   63949: out<=1;
   63950: out<=0;
   63951: out<=0;
   63952: out<=0;
   63953: out<=0;
   63954: out<=0;
   63955: out<=0;
   63956: out<=0;
   63957: out<=1;
   63958: out<=1;
   63959: out<=0;
   63960: out<=1;
   63961: out<=0;
   63962: out<=1;
   63963: out<=0;
   63964: out<=1;
   63965: out<=1;
   63966: out<=0;
   63967: out<=0;
   63968: out<=0;
   63969: out<=0;
   63970: out<=0;
   63971: out<=0;
   63972: out<=0;
   63973: out<=1;
   63974: out<=1;
   63975: out<=0;
   63976: out<=1;
   63977: out<=0;
   63978: out<=1;
   63979: out<=0;
   63980: out<=1;
   63981: out<=1;
   63982: out<=0;
   63983: out<=0;
   63984: out<=0;
   63985: out<=0;
   63986: out<=0;
   63987: out<=0;
   63988: out<=0;
   63989: out<=1;
   63990: out<=1;
   63991: out<=0;
   63992: out<=1;
   63993: out<=0;
   63994: out<=1;
   63995: out<=0;
   63996: out<=1;
   63997: out<=1;
   63998: out<=0;
   63999: out<=0;
   64000: out<=1;
   64001: out<=1;
   64002: out<=0;
   64003: out<=0;
   64004: out<=1;
   64005: out<=0;
   64006: out<=1;
   64007: out<=0;
   64008: out<=1;
   64009: out<=0;
   64010: out<=0;
   64011: out<=1;
   64012: out<=1;
   64013: out<=1;
   64014: out<=1;
   64015: out<=1;
   64016: out<=1;
   64017: out<=1;
   64018: out<=0;
   64019: out<=0;
   64020: out<=1;
   64021: out<=0;
   64022: out<=1;
   64023: out<=0;
   64024: out<=1;
   64025: out<=0;
   64026: out<=0;
   64027: out<=1;
   64028: out<=1;
   64029: out<=1;
   64030: out<=1;
   64031: out<=1;
   64032: out<=1;
   64033: out<=1;
   64034: out<=0;
   64035: out<=0;
   64036: out<=1;
   64037: out<=0;
   64038: out<=1;
   64039: out<=0;
   64040: out<=1;
   64041: out<=0;
   64042: out<=0;
   64043: out<=1;
   64044: out<=1;
   64045: out<=1;
   64046: out<=1;
   64047: out<=1;
   64048: out<=1;
   64049: out<=1;
   64050: out<=0;
   64051: out<=0;
   64052: out<=1;
   64053: out<=0;
   64054: out<=1;
   64055: out<=0;
   64056: out<=1;
   64057: out<=0;
   64058: out<=0;
   64059: out<=1;
   64060: out<=1;
   64061: out<=1;
   64062: out<=1;
   64063: out<=1;
   64064: out<=0;
   64065: out<=0;
   64066: out<=1;
   64067: out<=1;
   64068: out<=0;
   64069: out<=1;
   64070: out<=0;
   64071: out<=1;
   64072: out<=0;
   64073: out<=1;
   64074: out<=1;
   64075: out<=0;
   64076: out<=0;
   64077: out<=0;
   64078: out<=0;
   64079: out<=0;
   64080: out<=1;
   64081: out<=1;
   64082: out<=0;
   64083: out<=0;
   64084: out<=1;
   64085: out<=0;
   64086: out<=1;
   64087: out<=0;
   64088: out<=1;
   64089: out<=0;
   64090: out<=0;
   64091: out<=1;
   64092: out<=1;
   64093: out<=1;
   64094: out<=1;
   64095: out<=1;
   64096: out<=1;
   64097: out<=1;
   64098: out<=0;
   64099: out<=0;
   64100: out<=1;
   64101: out<=0;
   64102: out<=1;
   64103: out<=0;
   64104: out<=1;
   64105: out<=0;
   64106: out<=0;
   64107: out<=1;
   64108: out<=1;
   64109: out<=1;
   64110: out<=1;
   64111: out<=1;
   64112: out<=0;
   64113: out<=0;
   64114: out<=1;
   64115: out<=1;
   64116: out<=0;
   64117: out<=1;
   64118: out<=0;
   64119: out<=1;
   64120: out<=0;
   64121: out<=1;
   64122: out<=1;
   64123: out<=0;
   64124: out<=0;
   64125: out<=0;
   64126: out<=0;
   64127: out<=0;
   64128: out<=0;
   64129: out<=0;
   64130: out<=1;
   64131: out<=1;
   64132: out<=0;
   64133: out<=1;
   64134: out<=0;
   64135: out<=1;
   64136: out<=0;
   64137: out<=1;
   64138: out<=1;
   64139: out<=0;
   64140: out<=0;
   64141: out<=0;
   64142: out<=0;
   64143: out<=0;
   64144: out<=1;
   64145: out<=1;
   64146: out<=0;
   64147: out<=0;
   64148: out<=1;
   64149: out<=0;
   64150: out<=1;
   64151: out<=0;
   64152: out<=1;
   64153: out<=0;
   64154: out<=0;
   64155: out<=1;
   64156: out<=1;
   64157: out<=1;
   64158: out<=1;
   64159: out<=1;
   64160: out<=0;
   64161: out<=0;
   64162: out<=1;
   64163: out<=1;
   64164: out<=0;
   64165: out<=1;
   64166: out<=0;
   64167: out<=1;
   64168: out<=0;
   64169: out<=1;
   64170: out<=1;
   64171: out<=0;
   64172: out<=0;
   64173: out<=0;
   64174: out<=0;
   64175: out<=0;
   64176: out<=1;
   64177: out<=1;
   64178: out<=0;
   64179: out<=0;
   64180: out<=1;
   64181: out<=0;
   64182: out<=1;
   64183: out<=0;
   64184: out<=1;
   64185: out<=0;
   64186: out<=0;
   64187: out<=1;
   64188: out<=1;
   64189: out<=1;
   64190: out<=1;
   64191: out<=1;
   64192: out<=1;
   64193: out<=1;
   64194: out<=0;
   64195: out<=0;
   64196: out<=1;
   64197: out<=0;
   64198: out<=1;
   64199: out<=0;
   64200: out<=1;
   64201: out<=0;
   64202: out<=0;
   64203: out<=1;
   64204: out<=1;
   64205: out<=1;
   64206: out<=1;
   64207: out<=1;
   64208: out<=1;
   64209: out<=1;
   64210: out<=0;
   64211: out<=0;
   64212: out<=1;
   64213: out<=0;
   64214: out<=1;
   64215: out<=0;
   64216: out<=1;
   64217: out<=0;
   64218: out<=0;
   64219: out<=1;
   64220: out<=1;
   64221: out<=1;
   64222: out<=1;
   64223: out<=1;
   64224: out<=0;
   64225: out<=0;
   64226: out<=1;
   64227: out<=1;
   64228: out<=0;
   64229: out<=1;
   64230: out<=0;
   64231: out<=1;
   64232: out<=0;
   64233: out<=1;
   64234: out<=1;
   64235: out<=0;
   64236: out<=0;
   64237: out<=0;
   64238: out<=0;
   64239: out<=0;
   64240: out<=0;
   64241: out<=0;
   64242: out<=1;
   64243: out<=1;
   64244: out<=0;
   64245: out<=1;
   64246: out<=0;
   64247: out<=1;
   64248: out<=0;
   64249: out<=1;
   64250: out<=1;
   64251: out<=0;
   64252: out<=0;
   64253: out<=0;
   64254: out<=0;
   64255: out<=0;
   64256: out<=0;
   64257: out<=1;
   64258: out<=0;
   64259: out<=1;
   64260: out<=1;
   64261: out<=1;
   64262: out<=0;
   64263: out<=0;
   64264: out<=1;
   64265: out<=1;
   64266: out<=1;
   64267: out<=1;
   64268: out<=0;
   64269: out<=1;
   64270: out<=1;
   64271: out<=0;
   64272: out<=1;
   64273: out<=0;
   64274: out<=1;
   64275: out<=0;
   64276: out<=0;
   64277: out<=0;
   64278: out<=1;
   64279: out<=1;
   64280: out<=0;
   64281: out<=0;
   64282: out<=0;
   64283: out<=0;
   64284: out<=1;
   64285: out<=0;
   64286: out<=0;
   64287: out<=1;
   64288: out<=1;
   64289: out<=0;
   64290: out<=1;
   64291: out<=0;
   64292: out<=0;
   64293: out<=0;
   64294: out<=1;
   64295: out<=1;
   64296: out<=0;
   64297: out<=0;
   64298: out<=0;
   64299: out<=0;
   64300: out<=1;
   64301: out<=0;
   64302: out<=0;
   64303: out<=1;
   64304: out<=0;
   64305: out<=1;
   64306: out<=0;
   64307: out<=1;
   64308: out<=1;
   64309: out<=1;
   64310: out<=0;
   64311: out<=0;
   64312: out<=1;
   64313: out<=1;
   64314: out<=1;
   64315: out<=1;
   64316: out<=0;
   64317: out<=1;
   64318: out<=1;
   64319: out<=0;
   64320: out<=1;
   64321: out<=0;
   64322: out<=1;
   64323: out<=0;
   64324: out<=0;
   64325: out<=0;
   64326: out<=1;
   64327: out<=1;
   64328: out<=0;
   64329: out<=0;
   64330: out<=0;
   64331: out<=0;
   64332: out<=1;
   64333: out<=0;
   64334: out<=0;
   64335: out<=1;
   64336: out<=1;
   64337: out<=0;
   64338: out<=1;
   64339: out<=0;
   64340: out<=0;
   64341: out<=0;
   64342: out<=1;
   64343: out<=1;
   64344: out<=0;
   64345: out<=0;
   64346: out<=0;
   64347: out<=0;
   64348: out<=1;
   64349: out<=0;
   64350: out<=0;
   64351: out<=1;
   64352: out<=1;
   64353: out<=0;
   64354: out<=1;
   64355: out<=0;
   64356: out<=0;
   64357: out<=0;
   64358: out<=1;
   64359: out<=1;
   64360: out<=0;
   64361: out<=0;
   64362: out<=0;
   64363: out<=0;
   64364: out<=1;
   64365: out<=0;
   64366: out<=0;
   64367: out<=1;
   64368: out<=1;
   64369: out<=0;
   64370: out<=1;
   64371: out<=0;
   64372: out<=0;
   64373: out<=0;
   64374: out<=1;
   64375: out<=1;
   64376: out<=0;
   64377: out<=0;
   64378: out<=0;
   64379: out<=0;
   64380: out<=1;
   64381: out<=0;
   64382: out<=0;
   64383: out<=1;
   64384: out<=1;
   64385: out<=0;
   64386: out<=1;
   64387: out<=0;
   64388: out<=0;
   64389: out<=0;
   64390: out<=1;
   64391: out<=1;
   64392: out<=0;
   64393: out<=0;
   64394: out<=0;
   64395: out<=0;
   64396: out<=1;
   64397: out<=0;
   64398: out<=0;
   64399: out<=1;
   64400: out<=1;
   64401: out<=0;
   64402: out<=1;
   64403: out<=0;
   64404: out<=0;
   64405: out<=0;
   64406: out<=1;
   64407: out<=1;
   64408: out<=0;
   64409: out<=0;
   64410: out<=0;
   64411: out<=0;
   64412: out<=1;
   64413: out<=0;
   64414: out<=0;
   64415: out<=1;
   64416: out<=0;
   64417: out<=1;
   64418: out<=0;
   64419: out<=1;
   64420: out<=1;
   64421: out<=1;
   64422: out<=0;
   64423: out<=0;
   64424: out<=1;
   64425: out<=1;
   64426: out<=1;
   64427: out<=1;
   64428: out<=0;
   64429: out<=1;
   64430: out<=1;
   64431: out<=0;
   64432: out<=0;
   64433: out<=1;
   64434: out<=0;
   64435: out<=1;
   64436: out<=1;
   64437: out<=1;
   64438: out<=0;
   64439: out<=0;
   64440: out<=1;
   64441: out<=1;
   64442: out<=1;
   64443: out<=1;
   64444: out<=0;
   64445: out<=1;
   64446: out<=1;
   64447: out<=0;
   64448: out<=0;
   64449: out<=1;
   64450: out<=0;
   64451: out<=1;
   64452: out<=1;
   64453: out<=1;
   64454: out<=0;
   64455: out<=0;
   64456: out<=1;
   64457: out<=1;
   64458: out<=1;
   64459: out<=1;
   64460: out<=0;
   64461: out<=1;
   64462: out<=1;
   64463: out<=0;
   64464: out<=1;
   64465: out<=0;
   64466: out<=1;
   64467: out<=0;
   64468: out<=0;
   64469: out<=0;
   64470: out<=1;
   64471: out<=1;
   64472: out<=0;
   64473: out<=0;
   64474: out<=0;
   64475: out<=0;
   64476: out<=1;
   64477: out<=0;
   64478: out<=0;
   64479: out<=1;
   64480: out<=0;
   64481: out<=1;
   64482: out<=0;
   64483: out<=1;
   64484: out<=1;
   64485: out<=1;
   64486: out<=0;
   64487: out<=0;
   64488: out<=1;
   64489: out<=1;
   64490: out<=1;
   64491: out<=1;
   64492: out<=0;
   64493: out<=1;
   64494: out<=1;
   64495: out<=0;
   64496: out<=1;
   64497: out<=0;
   64498: out<=1;
   64499: out<=0;
   64500: out<=0;
   64501: out<=0;
   64502: out<=1;
   64503: out<=1;
   64504: out<=0;
   64505: out<=0;
   64506: out<=0;
   64507: out<=0;
   64508: out<=1;
   64509: out<=0;
   64510: out<=0;
   64511: out<=1;
   64512: out<=1;
   64513: out<=1;
   64514: out<=1;
   64515: out<=1;
   64516: out<=0;
   64517: out<=1;
   64518: out<=1;
   64519: out<=0;
   64520: out<=1;
   64521: out<=0;
   64522: out<=1;
   64523: out<=0;
   64524: out<=0;
   64525: out<=0;
   64526: out<=1;
   64527: out<=1;
   64528: out<=0;
   64529: out<=0;
   64530: out<=0;
   64531: out<=0;
   64532: out<=1;
   64533: out<=0;
   64534: out<=0;
   64535: out<=1;
   64536: out<=0;
   64537: out<=1;
   64538: out<=0;
   64539: out<=1;
   64540: out<=1;
   64541: out<=1;
   64542: out<=0;
   64543: out<=0;
   64544: out<=1;
   64545: out<=1;
   64546: out<=1;
   64547: out<=1;
   64548: out<=0;
   64549: out<=1;
   64550: out<=1;
   64551: out<=0;
   64552: out<=1;
   64553: out<=0;
   64554: out<=1;
   64555: out<=0;
   64556: out<=0;
   64557: out<=0;
   64558: out<=1;
   64559: out<=1;
   64560: out<=0;
   64561: out<=0;
   64562: out<=0;
   64563: out<=0;
   64564: out<=1;
   64565: out<=0;
   64566: out<=0;
   64567: out<=1;
   64568: out<=0;
   64569: out<=1;
   64570: out<=0;
   64571: out<=1;
   64572: out<=1;
   64573: out<=1;
   64574: out<=0;
   64575: out<=0;
   64576: out<=0;
   64577: out<=0;
   64578: out<=0;
   64579: out<=0;
   64580: out<=1;
   64581: out<=0;
   64582: out<=0;
   64583: out<=1;
   64584: out<=0;
   64585: out<=1;
   64586: out<=0;
   64587: out<=1;
   64588: out<=1;
   64589: out<=1;
   64590: out<=0;
   64591: out<=0;
   64592: out<=0;
   64593: out<=0;
   64594: out<=0;
   64595: out<=0;
   64596: out<=1;
   64597: out<=0;
   64598: out<=0;
   64599: out<=1;
   64600: out<=0;
   64601: out<=1;
   64602: out<=0;
   64603: out<=1;
   64604: out<=1;
   64605: out<=1;
   64606: out<=0;
   64607: out<=0;
   64608: out<=1;
   64609: out<=1;
   64610: out<=1;
   64611: out<=1;
   64612: out<=0;
   64613: out<=1;
   64614: out<=1;
   64615: out<=0;
   64616: out<=1;
   64617: out<=0;
   64618: out<=1;
   64619: out<=0;
   64620: out<=0;
   64621: out<=0;
   64622: out<=1;
   64623: out<=1;
   64624: out<=1;
   64625: out<=1;
   64626: out<=1;
   64627: out<=1;
   64628: out<=0;
   64629: out<=1;
   64630: out<=1;
   64631: out<=0;
   64632: out<=1;
   64633: out<=0;
   64634: out<=1;
   64635: out<=0;
   64636: out<=0;
   64637: out<=0;
   64638: out<=1;
   64639: out<=1;
   64640: out<=0;
   64641: out<=0;
   64642: out<=0;
   64643: out<=0;
   64644: out<=1;
   64645: out<=0;
   64646: out<=0;
   64647: out<=1;
   64648: out<=0;
   64649: out<=1;
   64650: out<=0;
   64651: out<=1;
   64652: out<=1;
   64653: out<=1;
   64654: out<=0;
   64655: out<=0;
   64656: out<=0;
   64657: out<=0;
   64658: out<=0;
   64659: out<=0;
   64660: out<=1;
   64661: out<=0;
   64662: out<=0;
   64663: out<=1;
   64664: out<=0;
   64665: out<=1;
   64666: out<=0;
   64667: out<=1;
   64668: out<=1;
   64669: out<=1;
   64670: out<=0;
   64671: out<=0;
   64672: out<=0;
   64673: out<=0;
   64674: out<=0;
   64675: out<=0;
   64676: out<=1;
   64677: out<=0;
   64678: out<=0;
   64679: out<=1;
   64680: out<=0;
   64681: out<=1;
   64682: out<=0;
   64683: out<=1;
   64684: out<=1;
   64685: out<=1;
   64686: out<=0;
   64687: out<=0;
   64688: out<=0;
   64689: out<=0;
   64690: out<=0;
   64691: out<=0;
   64692: out<=1;
   64693: out<=0;
   64694: out<=0;
   64695: out<=1;
   64696: out<=0;
   64697: out<=1;
   64698: out<=0;
   64699: out<=1;
   64700: out<=1;
   64701: out<=1;
   64702: out<=0;
   64703: out<=0;
   64704: out<=1;
   64705: out<=1;
   64706: out<=1;
   64707: out<=1;
   64708: out<=0;
   64709: out<=1;
   64710: out<=1;
   64711: out<=0;
   64712: out<=1;
   64713: out<=0;
   64714: out<=1;
   64715: out<=0;
   64716: out<=0;
   64717: out<=0;
   64718: out<=1;
   64719: out<=1;
   64720: out<=0;
   64721: out<=0;
   64722: out<=0;
   64723: out<=0;
   64724: out<=1;
   64725: out<=0;
   64726: out<=0;
   64727: out<=1;
   64728: out<=0;
   64729: out<=1;
   64730: out<=0;
   64731: out<=1;
   64732: out<=1;
   64733: out<=1;
   64734: out<=0;
   64735: out<=0;
   64736: out<=0;
   64737: out<=0;
   64738: out<=0;
   64739: out<=0;
   64740: out<=1;
   64741: out<=0;
   64742: out<=0;
   64743: out<=1;
   64744: out<=0;
   64745: out<=1;
   64746: out<=0;
   64747: out<=1;
   64748: out<=1;
   64749: out<=1;
   64750: out<=0;
   64751: out<=0;
   64752: out<=1;
   64753: out<=1;
   64754: out<=1;
   64755: out<=1;
   64756: out<=0;
   64757: out<=1;
   64758: out<=1;
   64759: out<=0;
   64760: out<=1;
   64761: out<=0;
   64762: out<=1;
   64763: out<=0;
   64764: out<=0;
   64765: out<=0;
   64766: out<=1;
   64767: out<=1;
   64768: out<=1;
   64769: out<=0;
   64770: out<=0;
   64771: out<=1;
   64772: out<=1;
   64773: out<=1;
   64774: out<=1;
   64775: out<=1;
   64776: out<=0;
   64777: out<=0;
   64778: out<=1;
   64779: out<=1;
   64780: out<=0;
   64781: out<=1;
   64782: out<=0;
   64783: out<=1;
   64784: out<=1;
   64785: out<=0;
   64786: out<=0;
   64787: out<=1;
   64788: out<=1;
   64789: out<=1;
   64790: out<=1;
   64791: out<=1;
   64792: out<=0;
   64793: out<=0;
   64794: out<=1;
   64795: out<=1;
   64796: out<=0;
   64797: out<=1;
   64798: out<=0;
   64799: out<=1;
   64800: out<=0;
   64801: out<=1;
   64802: out<=1;
   64803: out<=0;
   64804: out<=0;
   64805: out<=0;
   64806: out<=0;
   64807: out<=0;
   64808: out<=1;
   64809: out<=1;
   64810: out<=0;
   64811: out<=0;
   64812: out<=1;
   64813: out<=0;
   64814: out<=1;
   64815: out<=0;
   64816: out<=0;
   64817: out<=1;
   64818: out<=1;
   64819: out<=0;
   64820: out<=0;
   64821: out<=0;
   64822: out<=0;
   64823: out<=0;
   64824: out<=1;
   64825: out<=1;
   64826: out<=0;
   64827: out<=0;
   64828: out<=1;
   64829: out<=0;
   64830: out<=1;
   64831: out<=0;
   64832: out<=0;
   64833: out<=1;
   64834: out<=1;
   64835: out<=0;
   64836: out<=0;
   64837: out<=0;
   64838: out<=0;
   64839: out<=0;
   64840: out<=1;
   64841: out<=1;
   64842: out<=0;
   64843: out<=0;
   64844: out<=1;
   64845: out<=0;
   64846: out<=1;
   64847: out<=0;
   64848: out<=1;
   64849: out<=0;
   64850: out<=0;
   64851: out<=1;
   64852: out<=1;
   64853: out<=1;
   64854: out<=1;
   64855: out<=1;
   64856: out<=0;
   64857: out<=0;
   64858: out<=1;
   64859: out<=1;
   64860: out<=0;
   64861: out<=1;
   64862: out<=0;
   64863: out<=1;
   64864: out<=0;
   64865: out<=1;
   64866: out<=1;
   64867: out<=0;
   64868: out<=0;
   64869: out<=0;
   64870: out<=0;
   64871: out<=0;
   64872: out<=1;
   64873: out<=1;
   64874: out<=0;
   64875: out<=0;
   64876: out<=1;
   64877: out<=0;
   64878: out<=1;
   64879: out<=0;
   64880: out<=1;
   64881: out<=0;
   64882: out<=0;
   64883: out<=1;
   64884: out<=1;
   64885: out<=1;
   64886: out<=1;
   64887: out<=1;
   64888: out<=0;
   64889: out<=0;
   64890: out<=1;
   64891: out<=1;
   64892: out<=0;
   64893: out<=1;
   64894: out<=0;
   64895: out<=1;
   64896: out<=0;
   64897: out<=1;
   64898: out<=1;
   64899: out<=0;
   64900: out<=0;
   64901: out<=0;
   64902: out<=0;
   64903: out<=0;
   64904: out<=1;
   64905: out<=1;
   64906: out<=0;
   64907: out<=0;
   64908: out<=1;
   64909: out<=0;
   64910: out<=1;
   64911: out<=0;
   64912: out<=1;
   64913: out<=0;
   64914: out<=0;
   64915: out<=1;
   64916: out<=1;
   64917: out<=1;
   64918: out<=1;
   64919: out<=1;
   64920: out<=0;
   64921: out<=0;
   64922: out<=1;
   64923: out<=1;
   64924: out<=0;
   64925: out<=1;
   64926: out<=0;
   64927: out<=1;
   64928: out<=1;
   64929: out<=0;
   64930: out<=0;
   64931: out<=1;
   64932: out<=1;
   64933: out<=1;
   64934: out<=1;
   64935: out<=1;
   64936: out<=0;
   64937: out<=0;
   64938: out<=1;
   64939: out<=1;
   64940: out<=0;
   64941: out<=1;
   64942: out<=0;
   64943: out<=1;
   64944: out<=0;
   64945: out<=1;
   64946: out<=1;
   64947: out<=0;
   64948: out<=0;
   64949: out<=0;
   64950: out<=0;
   64951: out<=0;
   64952: out<=1;
   64953: out<=1;
   64954: out<=0;
   64955: out<=0;
   64956: out<=1;
   64957: out<=0;
   64958: out<=1;
   64959: out<=0;
   64960: out<=1;
   64961: out<=0;
   64962: out<=0;
   64963: out<=1;
   64964: out<=1;
   64965: out<=1;
   64966: out<=1;
   64967: out<=1;
   64968: out<=0;
   64969: out<=0;
   64970: out<=1;
   64971: out<=1;
   64972: out<=0;
   64973: out<=1;
   64974: out<=0;
   64975: out<=1;
   64976: out<=1;
   64977: out<=0;
   64978: out<=0;
   64979: out<=1;
   64980: out<=1;
   64981: out<=1;
   64982: out<=1;
   64983: out<=1;
   64984: out<=0;
   64985: out<=0;
   64986: out<=1;
   64987: out<=1;
   64988: out<=0;
   64989: out<=1;
   64990: out<=0;
   64991: out<=1;
   64992: out<=1;
   64993: out<=0;
   64994: out<=0;
   64995: out<=1;
   64996: out<=1;
   64997: out<=1;
   64998: out<=1;
   64999: out<=1;
   65000: out<=0;
   65001: out<=0;
   65002: out<=1;
   65003: out<=1;
   65004: out<=0;
   65005: out<=1;
   65006: out<=0;
   65007: out<=1;
   65008: out<=1;
   65009: out<=0;
   65010: out<=0;
   65011: out<=1;
   65012: out<=1;
   65013: out<=1;
   65014: out<=1;
   65015: out<=1;
   65016: out<=0;
   65017: out<=0;
   65018: out<=1;
   65019: out<=1;
   65020: out<=0;
   65021: out<=1;
   65022: out<=0;
   65023: out<=1;
   65024: out<=0;
   65025: out<=1;
   65026: out<=0;
   65027: out<=1;
   65028: out<=0;
   65029: out<=0;
   65030: out<=1;
   65031: out<=1;
   65032: out<=0;
   65033: out<=0;
   65034: out<=0;
   65035: out<=0;
   65036: out<=0;
   65037: out<=1;
   65038: out<=1;
   65039: out<=0;
   65040: out<=0;
   65041: out<=1;
   65042: out<=0;
   65043: out<=1;
   65044: out<=0;
   65045: out<=0;
   65046: out<=1;
   65047: out<=1;
   65048: out<=0;
   65049: out<=0;
   65050: out<=0;
   65051: out<=0;
   65052: out<=0;
   65053: out<=1;
   65054: out<=1;
   65055: out<=0;
   65056: out<=0;
   65057: out<=1;
   65058: out<=0;
   65059: out<=1;
   65060: out<=0;
   65061: out<=0;
   65062: out<=1;
   65063: out<=1;
   65064: out<=0;
   65065: out<=0;
   65066: out<=0;
   65067: out<=0;
   65068: out<=0;
   65069: out<=1;
   65070: out<=1;
   65071: out<=0;
   65072: out<=0;
   65073: out<=1;
   65074: out<=0;
   65075: out<=1;
   65076: out<=0;
   65077: out<=0;
   65078: out<=1;
   65079: out<=1;
   65080: out<=0;
   65081: out<=0;
   65082: out<=0;
   65083: out<=0;
   65084: out<=0;
   65085: out<=1;
   65086: out<=1;
   65087: out<=0;
   65088: out<=1;
   65089: out<=0;
   65090: out<=1;
   65091: out<=0;
   65092: out<=1;
   65093: out<=1;
   65094: out<=0;
   65095: out<=0;
   65096: out<=1;
   65097: out<=1;
   65098: out<=1;
   65099: out<=1;
   65100: out<=1;
   65101: out<=0;
   65102: out<=0;
   65103: out<=1;
   65104: out<=0;
   65105: out<=1;
   65106: out<=0;
   65107: out<=1;
   65108: out<=0;
   65109: out<=0;
   65110: out<=1;
   65111: out<=1;
   65112: out<=0;
   65113: out<=0;
   65114: out<=0;
   65115: out<=0;
   65116: out<=0;
   65117: out<=1;
   65118: out<=1;
   65119: out<=0;
   65120: out<=0;
   65121: out<=1;
   65122: out<=0;
   65123: out<=1;
   65124: out<=0;
   65125: out<=0;
   65126: out<=1;
   65127: out<=1;
   65128: out<=0;
   65129: out<=0;
   65130: out<=0;
   65131: out<=0;
   65132: out<=0;
   65133: out<=1;
   65134: out<=1;
   65135: out<=0;
   65136: out<=1;
   65137: out<=0;
   65138: out<=1;
   65139: out<=0;
   65140: out<=1;
   65141: out<=1;
   65142: out<=0;
   65143: out<=0;
   65144: out<=1;
   65145: out<=1;
   65146: out<=1;
   65147: out<=1;
   65148: out<=1;
   65149: out<=0;
   65150: out<=0;
   65151: out<=1;
   65152: out<=1;
   65153: out<=0;
   65154: out<=1;
   65155: out<=0;
   65156: out<=1;
   65157: out<=1;
   65158: out<=0;
   65159: out<=0;
   65160: out<=1;
   65161: out<=1;
   65162: out<=1;
   65163: out<=1;
   65164: out<=1;
   65165: out<=0;
   65166: out<=0;
   65167: out<=1;
   65168: out<=0;
   65169: out<=1;
   65170: out<=0;
   65171: out<=1;
   65172: out<=0;
   65173: out<=0;
   65174: out<=1;
   65175: out<=1;
   65176: out<=0;
   65177: out<=0;
   65178: out<=0;
   65179: out<=0;
   65180: out<=0;
   65181: out<=1;
   65182: out<=1;
   65183: out<=0;
   65184: out<=1;
   65185: out<=0;
   65186: out<=1;
   65187: out<=0;
   65188: out<=1;
   65189: out<=1;
   65190: out<=0;
   65191: out<=0;
   65192: out<=1;
   65193: out<=1;
   65194: out<=1;
   65195: out<=1;
   65196: out<=1;
   65197: out<=0;
   65198: out<=0;
   65199: out<=1;
   65200: out<=0;
   65201: out<=1;
   65202: out<=0;
   65203: out<=1;
   65204: out<=0;
   65205: out<=0;
   65206: out<=1;
   65207: out<=1;
   65208: out<=0;
   65209: out<=0;
   65210: out<=0;
   65211: out<=0;
   65212: out<=0;
   65213: out<=1;
   65214: out<=1;
   65215: out<=0;
   65216: out<=0;
   65217: out<=1;
   65218: out<=0;
   65219: out<=1;
   65220: out<=0;
   65221: out<=0;
   65222: out<=1;
   65223: out<=1;
   65224: out<=0;
   65225: out<=0;
   65226: out<=0;
   65227: out<=0;
   65228: out<=0;
   65229: out<=1;
   65230: out<=1;
   65231: out<=0;
   65232: out<=0;
   65233: out<=1;
   65234: out<=0;
   65235: out<=1;
   65236: out<=0;
   65237: out<=0;
   65238: out<=1;
   65239: out<=1;
   65240: out<=0;
   65241: out<=0;
   65242: out<=0;
   65243: out<=0;
   65244: out<=0;
   65245: out<=1;
   65246: out<=1;
   65247: out<=0;
   65248: out<=1;
   65249: out<=0;
   65250: out<=1;
   65251: out<=0;
   65252: out<=1;
   65253: out<=1;
   65254: out<=0;
   65255: out<=0;
   65256: out<=1;
   65257: out<=1;
   65258: out<=1;
   65259: out<=1;
   65260: out<=1;
   65261: out<=0;
   65262: out<=0;
   65263: out<=1;
   65264: out<=1;
   65265: out<=0;
   65266: out<=1;
   65267: out<=0;
   65268: out<=1;
   65269: out<=1;
   65270: out<=0;
   65271: out<=0;
   65272: out<=1;
   65273: out<=1;
   65274: out<=1;
   65275: out<=1;
   65276: out<=1;
   65277: out<=0;
   65278: out<=0;
   65279: out<=1;
   65280: out<=0;
   65281: out<=0;
   65282: out<=1;
   65283: out<=1;
   65284: out<=1;
   65285: out<=0;
   65286: out<=1;
   65287: out<=0;
   65288: out<=1;
   65289: out<=0;
   65290: out<=0;
   65291: out<=1;
   65292: out<=0;
   65293: out<=0;
   65294: out<=0;
   65295: out<=0;
   65296: out<=1;
   65297: out<=1;
   65298: out<=0;
   65299: out<=0;
   65300: out<=0;
   65301: out<=1;
   65302: out<=0;
   65303: out<=1;
   65304: out<=0;
   65305: out<=1;
   65306: out<=1;
   65307: out<=0;
   65308: out<=1;
   65309: out<=1;
   65310: out<=1;
   65311: out<=1;
   65312: out<=1;
   65313: out<=1;
   65314: out<=0;
   65315: out<=0;
   65316: out<=0;
   65317: out<=1;
   65318: out<=0;
   65319: out<=1;
   65320: out<=0;
   65321: out<=1;
   65322: out<=1;
   65323: out<=0;
   65324: out<=1;
   65325: out<=1;
   65326: out<=1;
   65327: out<=1;
   65328: out<=0;
   65329: out<=0;
   65330: out<=1;
   65331: out<=1;
   65332: out<=1;
   65333: out<=0;
   65334: out<=1;
   65335: out<=0;
   65336: out<=1;
   65337: out<=0;
   65338: out<=0;
   65339: out<=1;
   65340: out<=0;
   65341: out<=0;
   65342: out<=0;
   65343: out<=0;
   65344: out<=1;
   65345: out<=1;
   65346: out<=0;
   65347: out<=0;
   65348: out<=0;
   65349: out<=1;
   65350: out<=0;
   65351: out<=1;
   65352: out<=0;
   65353: out<=1;
   65354: out<=1;
   65355: out<=0;
   65356: out<=1;
   65357: out<=1;
   65358: out<=1;
   65359: out<=1;
   65360: out<=1;
   65361: out<=1;
   65362: out<=0;
   65363: out<=0;
   65364: out<=0;
   65365: out<=1;
   65366: out<=0;
   65367: out<=1;
   65368: out<=0;
   65369: out<=1;
   65370: out<=1;
   65371: out<=0;
   65372: out<=1;
   65373: out<=1;
   65374: out<=1;
   65375: out<=1;
   65376: out<=1;
   65377: out<=1;
   65378: out<=0;
   65379: out<=0;
   65380: out<=0;
   65381: out<=1;
   65382: out<=0;
   65383: out<=1;
   65384: out<=0;
   65385: out<=1;
   65386: out<=1;
   65387: out<=0;
   65388: out<=1;
   65389: out<=1;
   65390: out<=1;
   65391: out<=1;
   65392: out<=1;
   65393: out<=1;
   65394: out<=0;
   65395: out<=0;
   65396: out<=0;
   65397: out<=1;
   65398: out<=0;
   65399: out<=1;
   65400: out<=0;
   65401: out<=1;
   65402: out<=1;
   65403: out<=0;
   65404: out<=1;
   65405: out<=1;
   65406: out<=1;
   65407: out<=1;
   65408: out<=1;
   65409: out<=1;
   65410: out<=0;
   65411: out<=0;
   65412: out<=0;
   65413: out<=1;
   65414: out<=0;
   65415: out<=1;
   65416: out<=0;
   65417: out<=1;
   65418: out<=1;
   65419: out<=0;
   65420: out<=1;
   65421: out<=1;
   65422: out<=1;
   65423: out<=1;
   65424: out<=1;
   65425: out<=1;
   65426: out<=0;
   65427: out<=0;
   65428: out<=0;
   65429: out<=1;
   65430: out<=0;
   65431: out<=1;
   65432: out<=0;
   65433: out<=1;
   65434: out<=1;
   65435: out<=0;
   65436: out<=1;
   65437: out<=1;
   65438: out<=1;
   65439: out<=1;
   65440: out<=0;
   65441: out<=0;
   65442: out<=1;
   65443: out<=1;
   65444: out<=1;
   65445: out<=0;
   65446: out<=1;
   65447: out<=0;
   65448: out<=1;
   65449: out<=0;
   65450: out<=0;
   65451: out<=1;
   65452: out<=0;
   65453: out<=0;
   65454: out<=0;
   65455: out<=0;
   65456: out<=0;
   65457: out<=0;
   65458: out<=1;
   65459: out<=1;
   65460: out<=1;
   65461: out<=0;
   65462: out<=1;
   65463: out<=0;
   65464: out<=1;
   65465: out<=0;
   65466: out<=0;
   65467: out<=1;
   65468: out<=0;
   65469: out<=0;
   65470: out<=0;
   65471: out<=0;
   65472: out<=0;
   65473: out<=0;
   65474: out<=1;
   65475: out<=1;
   65476: out<=1;
   65477: out<=0;
   65478: out<=1;
   65479: out<=0;
   65480: out<=1;
   65481: out<=0;
   65482: out<=0;
   65483: out<=1;
   65484: out<=0;
   65485: out<=0;
   65486: out<=0;
   65487: out<=0;
   65488: out<=1;
   65489: out<=1;
   65490: out<=0;
   65491: out<=0;
   65492: out<=0;
   65493: out<=1;
   65494: out<=0;
   65495: out<=1;
   65496: out<=0;
   65497: out<=1;
   65498: out<=1;
   65499: out<=0;
   65500: out<=1;
   65501: out<=1;
   65502: out<=1;
   65503: out<=1;
   65504: out<=0;
   65505: out<=0;
   65506: out<=1;
   65507: out<=1;
   65508: out<=1;
   65509: out<=0;
   65510: out<=1;
   65511: out<=0;
   65512: out<=1;
   65513: out<=0;
   65514: out<=0;
   65515: out<=1;
   65516: out<=0;
   65517: out<=0;
   65518: out<=0;
   65519: out<=0;
   65520: out<=1;
   65521: out<=1;
   65522: out<=0;
   65523: out<=0;
   65524: out<=0;
   65525: out<=1;
   65526: out<=0;
   65527: out<=1;
   65528: out<=0;
   65529: out<=1;
   65530: out<=1;
   65531: out<=0;
   65532: out<=1;
   65533: out<=1;
   65534: out<=1;
   65535: out<=1;
 endcase
end
endmodule
