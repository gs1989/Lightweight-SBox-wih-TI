module STI8_R6_21487436(in,out);
  input[15:0] in;
  output out;
  reg out;
  always@(in)
  begin
    case(in)
   0: out<=0;
   1: out<=1;
   2: out<=0;
   3: out<=1;
   4: out<=0;
   5: out<=0;
   6: out<=1;
   7: out<=1;
   8: out<=0;
   9: out<=0;
   10: out<=0;
   11: out<=0;
   12: out<=0;
   13: out<=1;
   14: out<=1;
   15: out<=0;
   16: out<=1;
   17: out<=1;
   18: out<=0;
   19: out<=0;
   20: out<=0;
   21: out<=1;
   22: out<=0;
   23: out<=1;
   24: out<=0;
   25: out<=1;
   26: out<=1;
   27: out<=0;
   28: out<=1;
   29: out<=1;
   30: out<=1;
   31: out<=1;
   32: out<=0;
   33: out<=0;
   34: out<=0;
   35: out<=0;
   36: out<=1;
   37: out<=0;
   38: out<=0;
   39: out<=1;
   40: out<=0;
   41: out<=1;
   42: out<=0;
   43: out<=1;
   44: out<=1;
   45: out<=1;
   46: out<=0;
   47: out<=0;
   48: out<=1;
   49: out<=0;
   50: out<=0;
   51: out<=1;
   52: out<=1;
   53: out<=1;
   54: out<=1;
   55: out<=1;
   56: out<=0;
   57: out<=0;
   58: out<=1;
   59: out<=1;
   60: out<=0;
   61: out<=1;
   62: out<=0;
   63: out<=1;
   64: out<=1;
   65: out<=0;
   66: out<=1;
   67: out<=0;
   68: out<=1;
   69: out<=1;
   70: out<=0;
   71: out<=0;
   72: out<=1;
   73: out<=1;
   74: out<=1;
   75: out<=1;
   76: out<=1;
   77: out<=0;
   78: out<=0;
   79: out<=1;
   80: out<=1;
   81: out<=1;
   82: out<=0;
   83: out<=0;
   84: out<=0;
   85: out<=1;
   86: out<=0;
   87: out<=1;
   88: out<=0;
   89: out<=1;
   90: out<=1;
   91: out<=0;
   92: out<=1;
   93: out<=1;
   94: out<=1;
   95: out<=1;
   96: out<=0;
   97: out<=0;
   98: out<=0;
   99: out<=0;
   100: out<=1;
   101: out<=0;
   102: out<=0;
   103: out<=1;
   104: out<=0;
   105: out<=1;
   106: out<=0;
   107: out<=1;
   108: out<=1;
   109: out<=1;
   110: out<=0;
   111: out<=0;
   112: out<=0;
   113: out<=1;
   114: out<=1;
   115: out<=0;
   116: out<=0;
   117: out<=0;
   118: out<=0;
   119: out<=0;
   120: out<=1;
   121: out<=1;
   122: out<=0;
   123: out<=0;
   124: out<=1;
   125: out<=0;
   126: out<=1;
   127: out<=0;
   128: out<=0;
   129: out<=1;
   130: out<=0;
   131: out<=1;
   132: out<=0;
   133: out<=0;
   134: out<=1;
   135: out<=1;
   136: out<=0;
   137: out<=0;
   138: out<=0;
   139: out<=0;
   140: out<=0;
   141: out<=1;
   142: out<=1;
   143: out<=0;
   144: out<=0;
   145: out<=0;
   146: out<=1;
   147: out<=1;
   148: out<=1;
   149: out<=0;
   150: out<=1;
   151: out<=0;
   152: out<=1;
   153: out<=0;
   154: out<=0;
   155: out<=1;
   156: out<=0;
   157: out<=0;
   158: out<=0;
   159: out<=0;
   160: out<=0;
   161: out<=0;
   162: out<=0;
   163: out<=0;
   164: out<=1;
   165: out<=0;
   166: out<=0;
   167: out<=1;
   168: out<=0;
   169: out<=1;
   170: out<=0;
   171: out<=1;
   172: out<=1;
   173: out<=1;
   174: out<=0;
   175: out<=0;
   176: out<=0;
   177: out<=1;
   178: out<=1;
   179: out<=0;
   180: out<=0;
   181: out<=0;
   182: out<=0;
   183: out<=0;
   184: out<=1;
   185: out<=1;
   186: out<=0;
   187: out<=0;
   188: out<=1;
   189: out<=0;
   190: out<=1;
   191: out<=0;
   192: out<=1;
   193: out<=0;
   194: out<=1;
   195: out<=0;
   196: out<=1;
   197: out<=1;
   198: out<=0;
   199: out<=0;
   200: out<=1;
   201: out<=1;
   202: out<=1;
   203: out<=1;
   204: out<=1;
   205: out<=0;
   206: out<=0;
   207: out<=1;
   208: out<=0;
   209: out<=0;
   210: out<=1;
   211: out<=1;
   212: out<=1;
   213: out<=0;
   214: out<=1;
   215: out<=0;
   216: out<=1;
   217: out<=0;
   218: out<=0;
   219: out<=1;
   220: out<=0;
   221: out<=0;
   222: out<=0;
   223: out<=0;
   224: out<=0;
   225: out<=0;
   226: out<=0;
   227: out<=0;
   228: out<=1;
   229: out<=0;
   230: out<=0;
   231: out<=1;
   232: out<=0;
   233: out<=1;
   234: out<=0;
   235: out<=1;
   236: out<=1;
   237: out<=1;
   238: out<=0;
   239: out<=0;
   240: out<=1;
   241: out<=0;
   242: out<=0;
   243: out<=1;
   244: out<=1;
   245: out<=1;
   246: out<=1;
   247: out<=1;
   248: out<=0;
   249: out<=0;
   250: out<=1;
   251: out<=1;
   252: out<=0;
   253: out<=1;
   254: out<=0;
   255: out<=1;
   256: out<=1;
   257: out<=1;
   258: out<=0;
   259: out<=0;
   260: out<=0;
   261: out<=1;
   262: out<=0;
   263: out<=1;
   264: out<=0;
   265: out<=1;
   266: out<=1;
   267: out<=0;
   268: out<=1;
   269: out<=1;
   270: out<=1;
   271: out<=1;
   272: out<=1;
   273: out<=0;
   274: out<=1;
   275: out<=0;
   276: out<=1;
   277: out<=1;
   278: out<=0;
   279: out<=0;
   280: out<=1;
   281: out<=1;
   282: out<=1;
   283: out<=1;
   284: out<=1;
   285: out<=0;
   286: out<=0;
   287: out<=1;
   288: out<=0;
   289: out<=1;
   290: out<=1;
   291: out<=0;
   292: out<=0;
   293: out<=0;
   294: out<=0;
   295: out<=0;
   296: out<=1;
   297: out<=1;
   298: out<=0;
   299: out<=0;
   300: out<=1;
   301: out<=0;
   302: out<=1;
   303: out<=0;
   304: out<=0;
   305: out<=0;
   306: out<=0;
   307: out<=0;
   308: out<=1;
   309: out<=0;
   310: out<=0;
   311: out<=1;
   312: out<=0;
   313: out<=1;
   314: out<=0;
   315: out<=1;
   316: out<=1;
   317: out<=1;
   318: out<=0;
   319: out<=0;
   320: out<=1;
   321: out<=1;
   322: out<=0;
   323: out<=0;
   324: out<=0;
   325: out<=1;
   326: out<=0;
   327: out<=1;
   328: out<=0;
   329: out<=1;
   330: out<=1;
   331: out<=0;
   332: out<=1;
   333: out<=1;
   334: out<=1;
   335: out<=1;
   336: out<=0;
   337: out<=1;
   338: out<=0;
   339: out<=1;
   340: out<=0;
   341: out<=0;
   342: out<=1;
   343: out<=1;
   344: out<=0;
   345: out<=0;
   346: out<=0;
   347: out<=0;
   348: out<=0;
   349: out<=1;
   350: out<=1;
   351: out<=0;
   352: out<=1;
   353: out<=0;
   354: out<=0;
   355: out<=1;
   356: out<=1;
   357: out<=1;
   358: out<=1;
   359: out<=1;
   360: out<=0;
   361: out<=0;
   362: out<=1;
   363: out<=1;
   364: out<=0;
   365: out<=1;
   366: out<=0;
   367: out<=1;
   368: out<=0;
   369: out<=0;
   370: out<=0;
   371: out<=0;
   372: out<=1;
   373: out<=0;
   374: out<=0;
   375: out<=1;
   376: out<=0;
   377: out<=1;
   378: out<=0;
   379: out<=1;
   380: out<=1;
   381: out<=1;
   382: out<=0;
   383: out<=0;
   384: out<=0;
   385: out<=0;
   386: out<=1;
   387: out<=1;
   388: out<=1;
   389: out<=0;
   390: out<=1;
   391: out<=0;
   392: out<=1;
   393: out<=0;
   394: out<=0;
   395: out<=1;
   396: out<=0;
   397: out<=0;
   398: out<=0;
   399: out<=0;
   400: out<=1;
   401: out<=0;
   402: out<=1;
   403: out<=0;
   404: out<=1;
   405: out<=1;
   406: out<=0;
   407: out<=0;
   408: out<=1;
   409: out<=1;
   410: out<=1;
   411: out<=1;
   412: out<=1;
   413: out<=0;
   414: out<=0;
   415: out<=1;
   416: out<=1;
   417: out<=0;
   418: out<=0;
   419: out<=1;
   420: out<=1;
   421: out<=1;
   422: out<=1;
   423: out<=1;
   424: out<=0;
   425: out<=0;
   426: out<=1;
   427: out<=1;
   428: out<=0;
   429: out<=1;
   430: out<=0;
   431: out<=1;
   432: out<=0;
   433: out<=0;
   434: out<=0;
   435: out<=0;
   436: out<=1;
   437: out<=0;
   438: out<=0;
   439: out<=1;
   440: out<=0;
   441: out<=1;
   442: out<=0;
   443: out<=1;
   444: out<=1;
   445: out<=1;
   446: out<=0;
   447: out<=0;
   448: out<=0;
   449: out<=0;
   450: out<=1;
   451: out<=1;
   452: out<=1;
   453: out<=0;
   454: out<=1;
   455: out<=0;
   456: out<=1;
   457: out<=0;
   458: out<=0;
   459: out<=1;
   460: out<=0;
   461: out<=0;
   462: out<=0;
   463: out<=0;
   464: out<=0;
   465: out<=1;
   466: out<=0;
   467: out<=1;
   468: out<=0;
   469: out<=0;
   470: out<=1;
   471: out<=1;
   472: out<=0;
   473: out<=0;
   474: out<=0;
   475: out<=0;
   476: out<=0;
   477: out<=1;
   478: out<=1;
   479: out<=0;
   480: out<=0;
   481: out<=1;
   482: out<=1;
   483: out<=0;
   484: out<=0;
   485: out<=0;
   486: out<=0;
   487: out<=0;
   488: out<=1;
   489: out<=1;
   490: out<=0;
   491: out<=0;
   492: out<=1;
   493: out<=0;
   494: out<=1;
   495: out<=0;
   496: out<=0;
   497: out<=0;
   498: out<=0;
   499: out<=0;
   500: out<=1;
   501: out<=0;
   502: out<=0;
   503: out<=1;
   504: out<=0;
   505: out<=1;
   506: out<=0;
   507: out<=1;
   508: out<=1;
   509: out<=1;
   510: out<=0;
   511: out<=0;
   512: out<=0;
   513: out<=0;
   514: out<=0;
   515: out<=0;
   516: out<=1;
   517: out<=0;
   518: out<=0;
   519: out<=1;
   520: out<=0;
   521: out<=1;
   522: out<=0;
   523: out<=1;
   524: out<=1;
   525: out<=1;
   526: out<=0;
   527: out<=0;
   528: out<=0;
   529: out<=1;
   530: out<=1;
   531: out<=0;
   532: out<=0;
   533: out<=0;
   534: out<=0;
   535: out<=0;
   536: out<=1;
   537: out<=1;
   538: out<=0;
   539: out<=0;
   540: out<=1;
   541: out<=0;
   542: out<=1;
   543: out<=0;
   544: out<=0;
   545: out<=1;
   546: out<=0;
   547: out<=1;
   548: out<=0;
   549: out<=0;
   550: out<=1;
   551: out<=1;
   552: out<=0;
   553: out<=0;
   554: out<=0;
   555: out<=0;
   556: out<=0;
   557: out<=1;
   558: out<=1;
   559: out<=0;
   560: out<=0;
   561: out<=0;
   562: out<=1;
   563: out<=1;
   564: out<=1;
   565: out<=0;
   566: out<=1;
   567: out<=0;
   568: out<=1;
   569: out<=0;
   570: out<=0;
   571: out<=1;
   572: out<=0;
   573: out<=0;
   574: out<=0;
   575: out<=0;
   576: out<=0;
   577: out<=0;
   578: out<=0;
   579: out<=0;
   580: out<=1;
   581: out<=0;
   582: out<=0;
   583: out<=1;
   584: out<=0;
   585: out<=1;
   586: out<=0;
   587: out<=1;
   588: out<=1;
   589: out<=1;
   590: out<=0;
   591: out<=0;
   592: out<=1;
   593: out<=0;
   594: out<=0;
   595: out<=1;
   596: out<=1;
   597: out<=1;
   598: out<=1;
   599: out<=1;
   600: out<=0;
   601: out<=0;
   602: out<=1;
   603: out<=1;
   604: out<=0;
   605: out<=1;
   606: out<=0;
   607: out<=1;
   608: out<=1;
   609: out<=0;
   610: out<=1;
   611: out<=0;
   612: out<=1;
   613: out<=1;
   614: out<=0;
   615: out<=0;
   616: out<=1;
   617: out<=1;
   618: out<=1;
   619: out<=1;
   620: out<=1;
   621: out<=0;
   622: out<=0;
   623: out<=1;
   624: out<=0;
   625: out<=0;
   626: out<=1;
   627: out<=1;
   628: out<=1;
   629: out<=0;
   630: out<=1;
   631: out<=0;
   632: out<=1;
   633: out<=0;
   634: out<=0;
   635: out<=1;
   636: out<=0;
   637: out<=0;
   638: out<=0;
   639: out<=0;
   640: out<=0;
   641: out<=0;
   642: out<=0;
   643: out<=0;
   644: out<=1;
   645: out<=0;
   646: out<=0;
   647: out<=1;
   648: out<=0;
   649: out<=1;
   650: out<=0;
   651: out<=1;
   652: out<=1;
   653: out<=1;
   654: out<=0;
   655: out<=0;
   656: out<=1;
   657: out<=0;
   658: out<=0;
   659: out<=1;
   660: out<=1;
   661: out<=1;
   662: out<=1;
   663: out<=1;
   664: out<=0;
   665: out<=0;
   666: out<=1;
   667: out<=1;
   668: out<=0;
   669: out<=1;
   670: out<=0;
   671: out<=1;
   672: out<=0;
   673: out<=1;
   674: out<=0;
   675: out<=1;
   676: out<=0;
   677: out<=0;
   678: out<=1;
   679: out<=1;
   680: out<=0;
   681: out<=0;
   682: out<=0;
   683: out<=0;
   684: out<=0;
   685: out<=1;
   686: out<=1;
   687: out<=0;
   688: out<=1;
   689: out<=1;
   690: out<=0;
   691: out<=0;
   692: out<=0;
   693: out<=1;
   694: out<=0;
   695: out<=1;
   696: out<=0;
   697: out<=1;
   698: out<=1;
   699: out<=0;
   700: out<=1;
   701: out<=1;
   702: out<=1;
   703: out<=1;
   704: out<=0;
   705: out<=0;
   706: out<=0;
   707: out<=0;
   708: out<=1;
   709: out<=0;
   710: out<=0;
   711: out<=1;
   712: out<=0;
   713: out<=1;
   714: out<=0;
   715: out<=1;
   716: out<=1;
   717: out<=1;
   718: out<=0;
   719: out<=0;
   720: out<=0;
   721: out<=1;
   722: out<=1;
   723: out<=0;
   724: out<=0;
   725: out<=0;
   726: out<=0;
   727: out<=0;
   728: out<=1;
   729: out<=1;
   730: out<=0;
   731: out<=0;
   732: out<=1;
   733: out<=0;
   734: out<=1;
   735: out<=0;
   736: out<=1;
   737: out<=0;
   738: out<=1;
   739: out<=0;
   740: out<=1;
   741: out<=1;
   742: out<=0;
   743: out<=0;
   744: out<=1;
   745: out<=1;
   746: out<=1;
   747: out<=1;
   748: out<=1;
   749: out<=0;
   750: out<=0;
   751: out<=1;
   752: out<=1;
   753: out<=1;
   754: out<=0;
   755: out<=0;
   756: out<=0;
   757: out<=1;
   758: out<=0;
   759: out<=1;
   760: out<=0;
   761: out<=1;
   762: out<=1;
   763: out<=0;
   764: out<=1;
   765: out<=1;
   766: out<=1;
   767: out<=1;
   768: out<=1;
   769: out<=0;
   770: out<=0;
   771: out<=1;
   772: out<=1;
   773: out<=1;
   774: out<=1;
   775: out<=1;
   776: out<=0;
   777: out<=0;
   778: out<=1;
   779: out<=1;
   780: out<=0;
   781: out<=1;
   782: out<=0;
   783: out<=1;
   784: out<=0;
   785: out<=0;
   786: out<=0;
   787: out<=0;
   788: out<=1;
   789: out<=0;
   790: out<=0;
   791: out<=1;
   792: out<=0;
   793: out<=1;
   794: out<=0;
   795: out<=1;
   796: out<=1;
   797: out<=1;
   798: out<=0;
   799: out<=0;
   800: out<=0;
   801: out<=0;
   802: out<=1;
   803: out<=1;
   804: out<=1;
   805: out<=0;
   806: out<=1;
   807: out<=0;
   808: out<=1;
   809: out<=0;
   810: out<=0;
   811: out<=1;
   812: out<=0;
   813: out<=0;
   814: out<=0;
   815: out<=0;
   816: out<=1;
   817: out<=0;
   818: out<=1;
   819: out<=0;
   820: out<=1;
   821: out<=1;
   822: out<=0;
   823: out<=0;
   824: out<=1;
   825: out<=1;
   826: out<=1;
   827: out<=1;
   828: out<=1;
   829: out<=0;
   830: out<=0;
   831: out<=1;
   832: out<=0;
   833: out<=1;
   834: out<=1;
   835: out<=0;
   836: out<=0;
   837: out<=0;
   838: out<=0;
   839: out<=0;
   840: out<=1;
   841: out<=1;
   842: out<=0;
   843: out<=0;
   844: out<=1;
   845: out<=0;
   846: out<=1;
   847: out<=0;
   848: out<=0;
   849: out<=0;
   850: out<=0;
   851: out<=0;
   852: out<=1;
   853: out<=0;
   854: out<=0;
   855: out<=1;
   856: out<=0;
   857: out<=1;
   858: out<=0;
   859: out<=1;
   860: out<=1;
   861: out<=1;
   862: out<=0;
   863: out<=0;
   864: out<=0;
   865: out<=0;
   866: out<=1;
   867: out<=1;
   868: out<=1;
   869: out<=0;
   870: out<=1;
   871: out<=0;
   872: out<=1;
   873: out<=0;
   874: out<=0;
   875: out<=1;
   876: out<=0;
   877: out<=0;
   878: out<=0;
   879: out<=0;
   880: out<=0;
   881: out<=1;
   882: out<=0;
   883: out<=1;
   884: out<=0;
   885: out<=0;
   886: out<=1;
   887: out<=1;
   888: out<=0;
   889: out<=0;
   890: out<=0;
   891: out<=0;
   892: out<=0;
   893: out<=1;
   894: out<=1;
   895: out<=0;
   896: out<=0;
   897: out<=1;
   898: out<=1;
   899: out<=0;
   900: out<=0;
   901: out<=0;
   902: out<=0;
   903: out<=0;
   904: out<=1;
   905: out<=1;
   906: out<=0;
   907: out<=0;
   908: out<=1;
   909: out<=0;
   910: out<=1;
   911: out<=0;
   912: out<=0;
   913: out<=0;
   914: out<=0;
   915: out<=0;
   916: out<=1;
   917: out<=0;
   918: out<=0;
   919: out<=1;
   920: out<=0;
   921: out<=1;
   922: out<=0;
   923: out<=1;
   924: out<=1;
   925: out<=1;
   926: out<=0;
   927: out<=0;
   928: out<=1;
   929: out<=1;
   930: out<=0;
   931: out<=0;
   932: out<=0;
   933: out<=1;
   934: out<=0;
   935: out<=1;
   936: out<=0;
   937: out<=1;
   938: out<=1;
   939: out<=0;
   940: out<=1;
   941: out<=1;
   942: out<=1;
   943: out<=1;
   944: out<=1;
   945: out<=0;
   946: out<=1;
   947: out<=0;
   948: out<=1;
   949: out<=1;
   950: out<=0;
   951: out<=0;
   952: out<=1;
   953: out<=1;
   954: out<=1;
   955: out<=1;
   956: out<=1;
   957: out<=0;
   958: out<=0;
   959: out<=1;
   960: out<=1;
   961: out<=0;
   962: out<=0;
   963: out<=1;
   964: out<=1;
   965: out<=1;
   966: out<=1;
   967: out<=1;
   968: out<=0;
   969: out<=0;
   970: out<=1;
   971: out<=1;
   972: out<=0;
   973: out<=1;
   974: out<=0;
   975: out<=1;
   976: out<=0;
   977: out<=0;
   978: out<=0;
   979: out<=0;
   980: out<=1;
   981: out<=0;
   982: out<=0;
   983: out<=1;
   984: out<=0;
   985: out<=1;
   986: out<=0;
   987: out<=1;
   988: out<=1;
   989: out<=1;
   990: out<=0;
   991: out<=0;
   992: out<=1;
   993: out<=1;
   994: out<=0;
   995: out<=0;
   996: out<=0;
   997: out<=1;
   998: out<=0;
   999: out<=1;
   1000: out<=0;
   1001: out<=1;
   1002: out<=1;
   1003: out<=0;
   1004: out<=1;
   1005: out<=1;
   1006: out<=1;
   1007: out<=1;
   1008: out<=0;
   1009: out<=1;
   1010: out<=0;
   1011: out<=1;
   1012: out<=0;
   1013: out<=0;
   1014: out<=1;
   1015: out<=1;
   1016: out<=0;
   1017: out<=0;
   1018: out<=0;
   1019: out<=0;
   1020: out<=0;
   1021: out<=1;
   1022: out<=1;
   1023: out<=0;
   1024: out<=1;
   1025: out<=1;
   1026: out<=0;
   1027: out<=0;
   1028: out<=1;
   1029: out<=0;
   1030: out<=1;
   1031: out<=0;
   1032: out<=1;
   1033: out<=0;
   1034: out<=0;
   1035: out<=1;
   1036: out<=1;
   1037: out<=1;
   1038: out<=1;
   1039: out<=1;
   1040: out<=0;
   1041: out<=1;
   1042: out<=0;
   1043: out<=1;
   1044: out<=1;
   1045: out<=1;
   1046: out<=0;
   1047: out<=0;
   1048: out<=1;
   1049: out<=1;
   1050: out<=1;
   1051: out<=1;
   1052: out<=0;
   1053: out<=1;
   1054: out<=1;
   1055: out<=0;
   1056: out<=1;
   1057: out<=0;
   1058: out<=0;
   1059: out<=1;
   1060: out<=0;
   1061: out<=0;
   1062: out<=0;
   1063: out<=0;
   1064: out<=1;
   1065: out<=1;
   1066: out<=0;
   1067: out<=0;
   1068: out<=0;
   1069: out<=1;
   1070: out<=0;
   1071: out<=1;
   1072: out<=0;
   1073: out<=0;
   1074: out<=0;
   1075: out<=0;
   1076: out<=0;
   1077: out<=1;
   1078: out<=1;
   1079: out<=0;
   1080: out<=1;
   1081: out<=0;
   1082: out<=1;
   1083: out<=0;
   1084: out<=1;
   1085: out<=1;
   1086: out<=0;
   1087: out<=0;
   1088: out<=1;
   1089: out<=1;
   1090: out<=0;
   1091: out<=0;
   1092: out<=1;
   1093: out<=0;
   1094: out<=1;
   1095: out<=0;
   1096: out<=1;
   1097: out<=0;
   1098: out<=0;
   1099: out<=1;
   1100: out<=1;
   1101: out<=1;
   1102: out<=1;
   1103: out<=1;
   1104: out<=1;
   1105: out<=0;
   1106: out<=1;
   1107: out<=0;
   1108: out<=0;
   1109: out<=0;
   1110: out<=1;
   1111: out<=1;
   1112: out<=0;
   1113: out<=0;
   1114: out<=0;
   1115: out<=0;
   1116: out<=1;
   1117: out<=0;
   1118: out<=0;
   1119: out<=1;
   1120: out<=0;
   1121: out<=1;
   1122: out<=1;
   1123: out<=0;
   1124: out<=1;
   1125: out<=1;
   1126: out<=1;
   1127: out<=1;
   1128: out<=0;
   1129: out<=0;
   1130: out<=1;
   1131: out<=1;
   1132: out<=1;
   1133: out<=0;
   1134: out<=1;
   1135: out<=0;
   1136: out<=0;
   1137: out<=0;
   1138: out<=0;
   1139: out<=0;
   1140: out<=0;
   1141: out<=1;
   1142: out<=1;
   1143: out<=0;
   1144: out<=1;
   1145: out<=0;
   1146: out<=1;
   1147: out<=0;
   1148: out<=1;
   1149: out<=1;
   1150: out<=0;
   1151: out<=0;
   1152: out<=0;
   1153: out<=0;
   1154: out<=1;
   1155: out<=1;
   1156: out<=0;
   1157: out<=1;
   1158: out<=0;
   1159: out<=1;
   1160: out<=0;
   1161: out<=1;
   1162: out<=1;
   1163: out<=0;
   1164: out<=0;
   1165: out<=0;
   1166: out<=0;
   1167: out<=0;
   1168: out<=0;
   1169: out<=1;
   1170: out<=0;
   1171: out<=1;
   1172: out<=1;
   1173: out<=1;
   1174: out<=0;
   1175: out<=0;
   1176: out<=1;
   1177: out<=1;
   1178: out<=1;
   1179: out<=1;
   1180: out<=0;
   1181: out<=1;
   1182: out<=1;
   1183: out<=0;
   1184: out<=0;
   1185: out<=1;
   1186: out<=1;
   1187: out<=0;
   1188: out<=1;
   1189: out<=1;
   1190: out<=1;
   1191: out<=1;
   1192: out<=0;
   1193: out<=0;
   1194: out<=1;
   1195: out<=1;
   1196: out<=1;
   1197: out<=0;
   1198: out<=1;
   1199: out<=0;
   1200: out<=0;
   1201: out<=0;
   1202: out<=0;
   1203: out<=0;
   1204: out<=0;
   1205: out<=1;
   1206: out<=1;
   1207: out<=0;
   1208: out<=1;
   1209: out<=0;
   1210: out<=1;
   1211: out<=0;
   1212: out<=1;
   1213: out<=1;
   1214: out<=0;
   1215: out<=0;
   1216: out<=0;
   1217: out<=0;
   1218: out<=1;
   1219: out<=1;
   1220: out<=0;
   1221: out<=1;
   1222: out<=0;
   1223: out<=1;
   1224: out<=0;
   1225: out<=1;
   1226: out<=1;
   1227: out<=0;
   1228: out<=0;
   1229: out<=0;
   1230: out<=0;
   1231: out<=0;
   1232: out<=1;
   1233: out<=0;
   1234: out<=1;
   1235: out<=0;
   1236: out<=0;
   1237: out<=0;
   1238: out<=1;
   1239: out<=1;
   1240: out<=0;
   1241: out<=0;
   1242: out<=0;
   1243: out<=0;
   1244: out<=1;
   1245: out<=0;
   1246: out<=0;
   1247: out<=1;
   1248: out<=1;
   1249: out<=0;
   1250: out<=0;
   1251: out<=1;
   1252: out<=0;
   1253: out<=0;
   1254: out<=0;
   1255: out<=0;
   1256: out<=1;
   1257: out<=1;
   1258: out<=0;
   1259: out<=0;
   1260: out<=0;
   1261: out<=1;
   1262: out<=0;
   1263: out<=1;
   1264: out<=0;
   1265: out<=0;
   1266: out<=0;
   1267: out<=0;
   1268: out<=0;
   1269: out<=1;
   1270: out<=1;
   1271: out<=0;
   1272: out<=1;
   1273: out<=0;
   1274: out<=1;
   1275: out<=0;
   1276: out<=1;
   1277: out<=1;
   1278: out<=0;
   1279: out<=0;
   1280: out<=1;
   1281: out<=0;
   1282: out<=1;
   1283: out<=0;
   1284: out<=0;
   1285: out<=0;
   1286: out<=1;
   1287: out<=1;
   1288: out<=0;
   1289: out<=0;
   1290: out<=0;
   1291: out<=0;
   1292: out<=1;
   1293: out<=0;
   1294: out<=0;
   1295: out<=1;
   1296: out<=1;
   1297: out<=1;
   1298: out<=0;
   1299: out<=0;
   1300: out<=1;
   1301: out<=0;
   1302: out<=1;
   1303: out<=0;
   1304: out<=1;
   1305: out<=0;
   1306: out<=0;
   1307: out<=1;
   1308: out<=1;
   1309: out<=1;
   1310: out<=1;
   1311: out<=1;
   1312: out<=0;
   1313: out<=0;
   1314: out<=0;
   1315: out<=0;
   1316: out<=0;
   1317: out<=1;
   1318: out<=1;
   1319: out<=0;
   1320: out<=1;
   1321: out<=0;
   1322: out<=1;
   1323: out<=0;
   1324: out<=1;
   1325: out<=1;
   1326: out<=0;
   1327: out<=0;
   1328: out<=0;
   1329: out<=1;
   1330: out<=1;
   1331: out<=0;
   1332: out<=1;
   1333: out<=1;
   1334: out<=1;
   1335: out<=1;
   1336: out<=0;
   1337: out<=0;
   1338: out<=1;
   1339: out<=1;
   1340: out<=1;
   1341: out<=0;
   1342: out<=1;
   1343: out<=0;
   1344: out<=0;
   1345: out<=1;
   1346: out<=0;
   1347: out<=1;
   1348: out<=1;
   1349: out<=1;
   1350: out<=0;
   1351: out<=0;
   1352: out<=1;
   1353: out<=1;
   1354: out<=1;
   1355: out<=1;
   1356: out<=0;
   1357: out<=1;
   1358: out<=1;
   1359: out<=0;
   1360: out<=1;
   1361: out<=1;
   1362: out<=0;
   1363: out<=0;
   1364: out<=1;
   1365: out<=0;
   1366: out<=1;
   1367: out<=0;
   1368: out<=1;
   1369: out<=0;
   1370: out<=0;
   1371: out<=1;
   1372: out<=1;
   1373: out<=1;
   1374: out<=1;
   1375: out<=1;
   1376: out<=0;
   1377: out<=0;
   1378: out<=0;
   1379: out<=0;
   1380: out<=0;
   1381: out<=1;
   1382: out<=1;
   1383: out<=0;
   1384: out<=1;
   1385: out<=0;
   1386: out<=1;
   1387: out<=0;
   1388: out<=1;
   1389: out<=1;
   1390: out<=0;
   1391: out<=0;
   1392: out<=1;
   1393: out<=0;
   1394: out<=0;
   1395: out<=1;
   1396: out<=0;
   1397: out<=0;
   1398: out<=0;
   1399: out<=0;
   1400: out<=1;
   1401: out<=1;
   1402: out<=0;
   1403: out<=0;
   1404: out<=0;
   1405: out<=1;
   1406: out<=0;
   1407: out<=1;
   1408: out<=1;
   1409: out<=0;
   1410: out<=1;
   1411: out<=0;
   1412: out<=0;
   1413: out<=0;
   1414: out<=1;
   1415: out<=1;
   1416: out<=0;
   1417: out<=0;
   1418: out<=0;
   1419: out<=0;
   1420: out<=1;
   1421: out<=0;
   1422: out<=0;
   1423: out<=1;
   1424: out<=0;
   1425: out<=0;
   1426: out<=1;
   1427: out<=1;
   1428: out<=0;
   1429: out<=1;
   1430: out<=0;
   1431: out<=1;
   1432: out<=0;
   1433: out<=1;
   1434: out<=1;
   1435: out<=0;
   1436: out<=0;
   1437: out<=0;
   1438: out<=0;
   1439: out<=0;
   1440: out<=0;
   1441: out<=0;
   1442: out<=0;
   1443: out<=0;
   1444: out<=0;
   1445: out<=1;
   1446: out<=1;
   1447: out<=0;
   1448: out<=1;
   1449: out<=0;
   1450: out<=1;
   1451: out<=0;
   1452: out<=1;
   1453: out<=1;
   1454: out<=0;
   1455: out<=0;
   1456: out<=1;
   1457: out<=0;
   1458: out<=0;
   1459: out<=1;
   1460: out<=0;
   1461: out<=0;
   1462: out<=0;
   1463: out<=0;
   1464: out<=1;
   1465: out<=1;
   1466: out<=0;
   1467: out<=0;
   1468: out<=0;
   1469: out<=1;
   1470: out<=0;
   1471: out<=1;
   1472: out<=0;
   1473: out<=1;
   1474: out<=0;
   1475: out<=1;
   1476: out<=1;
   1477: out<=1;
   1478: out<=0;
   1479: out<=0;
   1480: out<=1;
   1481: out<=1;
   1482: out<=1;
   1483: out<=1;
   1484: out<=0;
   1485: out<=1;
   1486: out<=1;
   1487: out<=0;
   1488: out<=0;
   1489: out<=0;
   1490: out<=1;
   1491: out<=1;
   1492: out<=0;
   1493: out<=1;
   1494: out<=0;
   1495: out<=1;
   1496: out<=0;
   1497: out<=1;
   1498: out<=1;
   1499: out<=0;
   1500: out<=0;
   1501: out<=0;
   1502: out<=0;
   1503: out<=0;
   1504: out<=0;
   1505: out<=0;
   1506: out<=0;
   1507: out<=0;
   1508: out<=0;
   1509: out<=1;
   1510: out<=1;
   1511: out<=0;
   1512: out<=1;
   1513: out<=0;
   1514: out<=1;
   1515: out<=0;
   1516: out<=1;
   1517: out<=1;
   1518: out<=0;
   1519: out<=0;
   1520: out<=0;
   1521: out<=1;
   1522: out<=1;
   1523: out<=0;
   1524: out<=1;
   1525: out<=1;
   1526: out<=1;
   1527: out<=1;
   1528: out<=0;
   1529: out<=0;
   1530: out<=1;
   1531: out<=1;
   1532: out<=1;
   1533: out<=0;
   1534: out<=1;
   1535: out<=0;
   1536: out<=0;
   1537: out<=1;
   1538: out<=1;
   1539: out<=0;
   1540: out<=1;
   1541: out<=1;
   1542: out<=1;
   1543: out<=1;
   1544: out<=0;
   1545: out<=0;
   1546: out<=1;
   1547: out<=1;
   1548: out<=1;
   1549: out<=0;
   1550: out<=1;
   1551: out<=0;
   1552: out<=0;
   1553: out<=0;
   1554: out<=0;
   1555: out<=0;
   1556: out<=0;
   1557: out<=1;
   1558: out<=1;
   1559: out<=0;
   1560: out<=1;
   1561: out<=0;
   1562: out<=1;
   1563: out<=0;
   1564: out<=1;
   1565: out<=1;
   1566: out<=0;
   1567: out<=0;
   1568: out<=0;
   1569: out<=0;
   1570: out<=1;
   1571: out<=1;
   1572: out<=0;
   1573: out<=1;
   1574: out<=0;
   1575: out<=1;
   1576: out<=0;
   1577: out<=1;
   1578: out<=1;
   1579: out<=0;
   1580: out<=0;
   1581: out<=0;
   1582: out<=0;
   1583: out<=0;
   1584: out<=0;
   1585: out<=1;
   1586: out<=0;
   1587: out<=1;
   1588: out<=1;
   1589: out<=1;
   1590: out<=0;
   1591: out<=0;
   1592: out<=1;
   1593: out<=1;
   1594: out<=1;
   1595: out<=1;
   1596: out<=0;
   1597: out<=1;
   1598: out<=1;
   1599: out<=0;
   1600: out<=1;
   1601: out<=0;
   1602: out<=0;
   1603: out<=1;
   1604: out<=0;
   1605: out<=0;
   1606: out<=0;
   1607: out<=0;
   1608: out<=1;
   1609: out<=1;
   1610: out<=0;
   1611: out<=0;
   1612: out<=0;
   1613: out<=1;
   1614: out<=0;
   1615: out<=1;
   1616: out<=0;
   1617: out<=0;
   1618: out<=0;
   1619: out<=0;
   1620: out<=0;
   1621: out<=1;
   1622: out<=1;
   1623: out<=0;
   1624: out<=1;
   1625: out<=0;
   1626: out<=1;
   1627: out<=0;
   1628: out<=1;
   1629: out<=1;
   1630: out<=0;
   1631: out<=0;
   1632: out<=0;
   1633: out<=0;
   1634: out<=1;
   1635: out<=1;
   1636: out<=0;
   1637: out<=1;
   1638: out<=0;
   1639: out<=1;
   1640: out<=0;
   1641: out<=1;
   1642: out<=1;
   1643: out<=0;
   1644: out<=0;
   1645: out<=0;
   1646: out<=0;
   1647: out<=0;
   1648: out<=1;
   1649: out<=0;
   1650: out<=1;
   1651: out<=0;
   1652: out<=0;
   1653: out<=0;
   1654: out<=1;
   1655: out<=1;
   1656: out<=0;
   1657: out<=0;
   1658: out<=0;
   1659: out<=0;
   1660: out<=1;
   1661: out<=0;
   1662: out<=0;
   1663: out<=1;
   1664: out<=1;
   1665: out<=0;
   1666: out<=0;
   1667: out<=1;
   1668: out<=0;
   1669: out<=0;
   1670: out<=0;
   1671: out<=0;
   1672: out<=1;
   1673: out<=1;
   1674: out<=0;
   1675: out<=0;
   1676: out<=0;
   1677: out<=1;
   1678: out<=0;
   1679: out<=1;
   1680: out<=0;
   1681: out<=0;
   1682: out<=0;
   1683: out<=0;
   1684: out<=0;
   1685: out<=1;
   1686: out<=1;
   1687: out<=0;
   1688: out<=1;
   1689: out<=0;
   1690: out<=1;
   1691: out<=0;
   1692: out<=1;
   1693: out<=1;
   1694: out<=0;
   1695: out<=0;
   1696: out<=1;
   1697: out<=1;
   1698: out<=0;
   1699: out<=0;
   1700: out<=1;
   1701: out<=0;
   1702: out<=1;
   1703: out<=0;
   1704: out<=1;
   1705: out<=0;
   1706: out<=0;
   1707: out<=1;
   1708: out<=1;
   1709: out<=1;
   1710: out<=1;
   1711: out<=1;
   1712: out<=0;
   1713: out<=1;
   1714: out<=0;
   1715: out<=1;
   1716: out<=1;
   1717: out<=1;
   1718: out<=0;
   1719: out<=0;
   1720: out<=1;
   1721: out<=1;
   1722: out<=1;
   1723: out<=1;
   1724: out<=0;
   1725: out<=1;
   1726: out<=1;
   1727: out<=0;
   1728: out<=0;
   1729: out<=1;
   1730: out<=1;
   1731: out<=0;
   1732: out<=1;
   1733: out<=1;
   1734: out<=1;
   1735: out<=1;
   1736: out<=0;
   1737: out<=0;
   1738: out<=1;
   1739: out<=1;
   1740: out<=1;
   1741: out<=0;
   1742: out<=1;
   1743: out<=0;
   1744: out<=0;
   1745: out<=0;
   1746: out<=0;
   1747: out<=0;
   1748: out<=0;
   1749: out<=1;
   1750: out<=1;
   1751: out<=0;
   1752: out<=1;
   1753: out<=0;
   1754: out<=1;
   1755: out<=0;
   1756: out<=1;
   1757: out<=1;
   1758: out<=0;
   1759: out<=0;
   1760: out<=1;
   1761: out<=1;
   1762: out<=0;
   1763: out<=0;
   1764: out<=1;
   1765: out<=0;
   1766: out<=1;
   1767: out<=0;
   1768: out<=1;
   1769: out<=0;
   1770: out<=0;
   1771: out<=1;
   1772: out<=1;
   1773: out<=1;
   1774: out<=1;
   1775: out<=1;
   1776: out<=1;
   1777: out<=0;
   1778: out<=1;
   1779: out<=0;
   1780: out<=0;
   1781: out<=0;
   1782: out<=1;
   1783: out<=1;
   1784: out<=0;
   1785: out<=0;
   1786: out<=0;
   1787: out<=0;
   1788: out<=1;
   1789: out<=0;
   1790: out<=0;
   1791: out<=1;
   1792: out<=0;
   1793: out<=0;
   1794: out<=0;
   1795: out<=0;
   1796: out<=0;
   1797: out<=1;
   1798: out<=1;
   1799: out<=0;
   1800: out<=1;
   1801: out<=0;
   1802: out<=1;
   1803: out<=0;
   1804: out<=1;
   1805: out<=1;
   1806: out<=0;
   1807: out<=0;
   1808: out<=1;
   1809: out<=0;
   1810: out<=0;
   1811: out<=1;
   1812: out<=0;
   1813: out<=0;
   1814: out<=0;
   1815: out<=0;
   1816: out<=1;
   1817: out<=1;
   1818: out<=0;
   1819: out<=0;
   1820: out<=0;
   1821: out<=1;
   1822: out<=0;
   1823: out<=1;
   1824: out<=1;
   1825: out<=0;
   1826: out<=1;
   1827: out<=0;
   1828: out<=0;
   1829: out<=0;
   1830: out<=1;
   1831: out<=1;
   1832: out<=0;
   1833: out<=0;
   1834: out<=0;
   1835: out<=0;
   1836: out<=1;
   1837: out<=0;
   1838: out<=0;
   1839: out<=1;
   1840: out<=0;
   1841: out<=0;
   1842: out<=1;
   1843: out<=1;
   1844: out<=0;
   1845: out<=1;
   1846: out<=0;
   1847: out<=1;
   1848: out<=0;
   1849: out<=1;
   1850: out<=1;
   1851: out<=0;
   1852: out<=0;
   1853: out<=0;
   1854: out<=0;
   1855: out<=0;
   1856: out<=0;
   1857: out<=0;
   1858: out<=0;
   1859: out<=0;
   1860: out<=0;
   1861: out<=1;
   1862: out<=1;
   1863: out<=0;
   1864: out<=1;
   1865: out<=0;
   1866: out<=1;
   1867: out<=0;
   1868: out<=1;
   1869: out<=1;
   1870: out<=0;
   1871: out<=0;
   1872: out<=0;
   1873: out<=1;
   1874: out<=1;
   1875: out<=0;
   1876: out<=1;
   1877: out<=1;
   1878: out<=1;
   1879: out<=1;
   1880: out<=0;
   1881: out<=0;
   1882: out<=1;
   1883: out<=1;
   1884: out<=1;
   1885: out<=0;
   1886: out<=1;
   1887: out<=0;
   1888: out<=0;
   1889: out<=1;
   1890: out<=0;
   1891: out<=1;
   1892: out<=1;
   1893: out<=1;
   1894: out<=0;
   1895: out<=0;
   1896: out<=1;
   1897: out<=1;
   1898: out<=1;
   1899: out<=1;
   1900: out<=0;
   1901: out<=1;
   1902: out<=1;
   1903: out<=0;
   1904: out<=0;
   1905: out<=0;
   1906: out<=1;
   1907: out<=1;
   1908: out<=0;
   1909: out<=1;
   1910: out<=0;
   1911: out<=1;
   1912: out<=0;
   1913: out<=1;
   1914: out<=1;
   1915: out<=0;
   1916: out<=0;
   1917: out<=0;
   1918: out<=0;
   1919: out<=0;
   1920: out<=0;
   1921: out<=0;
   1922: out<=0;
   1923: out<=0;
   1924: out<=0;
   1925: out<=1;
   1926: out<=1;
   1927: out<=0;
   1928: out<=1;
   1929: out<=0;
   1930: out<=1;
   1931: out<=0;
   1932: out<=1;
   1933: out<=1;
   1934: out<=0;
   1935: out<=0;
   1936: out<=0;
   1937: out<=1;
   1938: out<=1;
   1939: out<=0;
   1940: out<=1;
   1941: out<=1;
   1942: out<=1;
   1943: out<=1;
   1944: out<=0;
   1945: out<=0;
   1946: out<=1;
   1947: out<=1;
   1948: out<=1;
   1949: out<=0;
   1950: out<=1;
   1951: out<=0;
   1952: out<=1;
   1953: out<=0;
   1954: out<=1;
   1955: out<=0;
   1956: out<=0;
   1957: out<=0;
   1958: out<=1;
   1959: out<=1;
   1960: out<=0;
   1961: out<=0;
   1962: out<=0;
   1963: out<=0;
   1964: out<=1;
   1965: out<=0;
   1966: out<=0;
   1967: out<=1;
   1968: out<=1;
   1969: out<=1;
   1970: out<=0;
   1971: out<=0;
   1972: out<=1;
   1973: out<=0;
   1974: out<=1;
   1975: out<=0;
   1976: out<=1;
   1977: out<=0;
   1978: out<=0;
   1979: out<=1;
   1980: out<=1;
   1981: out<=1;
   1982: out<=1;
   1983: out<=1;
   1984: out<=0;
   1985: out<=0;
   1986: out<=0;
   1987: out<=0;
   1988: out<=0;
   1989: out<=1;
   1990: out<=1;
   1991: out<=0;
   1992: out<=1;
   1993: out<=0;
   1994: out<=1;
   1995: out<=0;
   1996: out<=1;
   1997: out<=1;
   1998: out<=0;
   1999: out<=0;
   2000: out<=1;
   2001: out<=0;
   2002: out<=0;
   2003: out<=1;
   2004: out<=0;
   2005: out<=0;
   2006: out<=0;
   2007: out<=0;
   2008: out<=1;
   2009: out<=1;
   2010: out<=0;
   2011: out<=0;
   2012: out<=0;
   2013: out<=1;
   2014: out<=0;
   2015: out<=1;
   2016: out<=0;
   2017: out<=1;
   2018: out<=0;
   2019: out<=1;
   2020: out<=1;
   2021: out<=1;
   2022: out<=0;
   2023: out<=0;
   2024: out<=1;
   2025: out<=1;
   2026: out<=1;
   2027: out<=1;
   2028: out<=0;
   2029: out<=1;
   2030: out<=1;
   2031: out<=0;
   2032: out<=1;
   2033: out<=1;
   2034: out<=0;
   2035: out<=0;
   2036: out<=1;
   2037: out<=0;
   2038: out<=1;
   2039: out<=0;
   2040: out<=1;
   2041: out<=0;
   2042: out<=0;
   2043: out<=1;
   2044: out<=1;
   2045: out<=1;
   2046: out<=1;
   2047: out<=1;
   2048: out<=0;
   2049: out<=0;
   2050: out<=0;
   2051: out<=0;
   2052: out<=0;
   2053: out<=1;
   2054: out<=1;
   2055: out<=0;
   2056: out<=0;
   2057: out<=1;
   2058: out<=0;
   2059: out<=1;
   2060: out<=0;
   2061: out<=0;
   2062: out<=1;
   2063: out<=1;
   2064: out<=1;
   2065: out<=0;
   2066: out<=0;
   2067: out<=1;
   2068: out<=0;
   2069: out<=0;
   2070: out<=0;
   2071: out<=0;
   2072: out<=0;
   2073: out<=0;
   2074: out<=1;
   2075: out<=1;
   2076: out<=1;
   2077: out<=0;
   2078: out<=1;
   2079: out<=0;
   2080: out<=0;
   2081: out<=1;
   2082: out<=0;
   2083: out<=1;
   2084: out<=1;
   2085: out<=1;
   2086: out<=0;
   2087: out<=0;
   2088: out<=0;
   2089: out<=0;
   2090: out<=0;
   2091: out<=0;
   2092: out<=1;
   2093: out<=0;
   2094: out<=0;
   2095: out<=1;
   2096: out<=1;
   2097: out<=1;
   2098: out<=0;
   2099: out<=0;
   2100: out<=1;
   2101: out<=0;
   2102: out<=1;
   2103: out<=0;
   2104: out<=0;
   2105: out<=1;
   2106: out<=1;
   2107: out<=0;
   2108: out<=0;
   2109: out<=0;
   2110: out<=0;
   2111: out<=0;
   2112: out<=0;
   2113: out<=0;
   2114: out<=0;
   2115: out<=0;
   2116: out<=0;
   2117: out<=1;
   2118: out<=1;
   2119: out<=0;
   2120: out<=0;
   2121: out<=1;
   2122: out<=0;
   2123: out<=1;
   2124: out<=0;
   2125: out<=0;
   2126: out<=1;
   2127: out<=1;
   2128: out<=0;
   2129: out<=1;
   2130: out<=1;
   2131: out<=0;
   2132: out<=1;
   2133: out<=1;
   2134: out<=1;
   2135: out<=1;
   2136: out<=1;
   2137: out<=1;
   2138: out<=0;
   2139: out<=0;
   2140: out<=0;
   2141: out<=1;
   2142: out<=0;
   2143: out<=1;
   2144: out<=1;
   2145: out<=0;
   2146: out<=1;
   2147: out<=0;
   2148: out<=0;
   2149: out<=0;
   2150: out<=1;
   2151: out<=1;
   2152: out<=1;
   2153: out<=1;
   2154: out<=1;
   2155: out<=1;
   2156: out<=0;
   2157: out<=1;
   2158: out<=1;
   2159: out<=0;
   2160: out<=1;
   2161: out<=1;
   2162: out<=0;
   2163: out<=0;
   2164: out<=1;
   2165: out<=0;
   2166: out<=1;
   2167: out<=0;
   2168: out<=0;
   2169: out<=1;
   2170: out<=1;
   2171: out<=0;
   2172: out<=0;
   2173: out<=0;
   2174: out<=0;
   2175: out<=0;
   2176: out<=0;
   2177: out<=0;
   2178: out<=0;
   2179: out<=0;
   2180: out<=0;
   2181: out<=1;
   2182: out<=1;
   2183: out<=0;
   2184: out<=0;
   2185: out<=1;
   2186: out<=0;
   2187: out<=1;
   2188: out<=0;
   2189: out<=0;
   2190: out<=1;
   2191: out<=1;
   2192: out<=0;
   2193: out<=1;
   2194: out<=1;
   2195: out<=0;
   2196: out<=1;
   2197: out<=1;
   2198: out<=1;
   2199: out<=1;
   2200: out<=1;
   2201: out<=1;
   2202: out<=0;
   2203: out<=0;
   2204: out<=0;
   2205: out<=1;
   2206: out<=0;
   2207: out<=1;
   2208: out<=0;
   2209: out<=1;
   2210: out<=0;
   2211: out<=1;
   2212: out<=1;
   2213: out<=1;
   2214: out<=0;
   2215: out<=0;
   2216: out<=0;
   2217: out<=0;
   2218: out<=0;
   2219: out<=0;
   2220: out<=1;
   2221: out<=0;
   2222: out<=0;
   2223: out<=1;
   2224: out<=0;
   2225: out<=0;
   2226: out<=1;
   2227: out<=1;
   2228: out<=0;
   2229: out<=1;
   2230: out<=0;
   2231: out<=1;
   2232: out<=1;
   2233: out<=0;
   2234: out<=0;
   2235: out<=1;
   2236: out<=1;
   2237: out<=1;
   2238: out<=1;
   2239: out<=1;
   2240: out<=0;
   2241: out<=0;
   2242: out<=0;
   2243: out<=0;
   2244: out<=0;
   2245: out<=1;
   2246: out<=1;
   2247: out<=0;
   2248: out<=0;
   2249: out<=1;
   2250: out<=0;
   2251: out<=1;
   2252: out<=0;
   2253: out<=0;
   2254: out<=1;
   2255: out<=1;
   2256: out<=1;
   2257: out<=0;
   2258: out<=0;
   2259: out<=1;
   2260: out<=0;
   2261: out<=0;
   2262: out<=0;
   2263: out<=0;
   2264: out<=0;
   2265: out<=0;
   2266: out<=1;
   2267: out<=1;
   2268: out<=1;
   2269: out<=0;
   2270: out<=1;
   2271: out<=0;
   2272: out<=1;
   2273: out<=0;
   2274: out<=1;
   2275: out<=0;
   2276: out<=0;
   2277: out<=0;
   2278: out<=1;
   2279: out<=1;
   2280: out<=1;
   2281: out<=1;
   2282: out<=1;
   2283: out<=1;
   2284: out<=0;
   2285: out<=1;
   2286: out<=1;
   2287: out<=0;
   2288: out<=0;
   2289: out<=0;
   2290: out<=1;
   2291: out<=1;
   2292: out<=0;
   2293: out<=1;
   2294: out<=0;
   2295: out<=1;
   2296: out<=1;
   2297: out<=0;
   2298: out<=0;
   2299: out<=1;
   2300: out<=1;
   2301: out<=1;
   2302: out<=1;
   2303: out<=1;
   2304: out<=0;
   2305: out<=1;
   2306: out<=1;
   2307: out<=0;
   2308: out<=1;
   2309: out<=1;
   2310: out<=1;
   2311: out<=1;
   2312: out<=1;
   2313: out<=1;
   2314: out<=0;
   2315: out<=0;
   2316: out<=0;
   2317: out<=1;
   2318: out<=0;
   2319: out<=1;
   2320: out<=0;
   2321: out<=0;
   2322: out<=0;
   2323: out<=0;
   2324: out<=0;
   2325: out<=1;
   2326: out<=1;
   2327: out<=0;
   2328: out<=0;
   2329: out<=1;
   2330: out<=0;
   2331: out<=1;
   2332: out<=0;
   2333: out<=0;
   2334: out<=1;
   2335: out<=1;
   2336: out<=1;
   2337: out<=1;
   2338: out<=0;
   2339: out<=0;
   2340: out<=1;
   2341: out<=0;
   2342: out<=1;
   2343: out<=0;
   2344: out<=0;
   2345: out<=1;
   2346: out<=1;
   2347: out<=0;
   2348: out<=0;
   2349: out<=0;
   2350: out<=0;
   2351: out<=0;
   2352: out<=1;
   2353: out<=0;
   2354: out<=1;
   2355: out<=0;
   2356: out<=0;
   2357: out<=0;
   2358: out<=1;
   2359: out<=1;
   2360: out<=1;
   2361: out<=1;
   2362: out<=1;
   2363: out<=1;
   2364: out<=0;
   2365: out<=1;
   2366: out<=1;
   2367: out<=0;
   2368: out<=1;
   2369: out<=0;
   2370: out<=0;
   2371: out<=1;
   2372: out<=0;
   2373: out<=0;
   2374: out<=0;
   2375: out<=0;
   2376: out<=0;
   2377: out<=0;
   2378: out<=1;
   2379: out<=1;
   2380: out<=1;
   2381: out<=0;
   2382: out<=1;
   2383: out<=0;
   2384: out<=0;
   2385: out<=0;
   2386: out<=0;
   2387: out<=0;
   2388: out<=0;
   2389: out<=1;
   2390: out<=1;
   2391: out<=0;
   2392: out<=0;
   2393: out<=1;
   2394: out<=0;
   2395: out<=1;
   2396: out<=0;
   2397: out<=0;
   2398: out<=1;
   2399: out<=1;
   2400: out<=1;
   2401: out<=1;
   2402: out<=0;
   2403: out<=0;
   2404: out<=1;
   2405: out<=0;
   2406: out<=1;
   2407: out<=0;
   2408: out<=0;
   2409: out<=1;
   2410: out<=1;
   2411: out<=0;
   2412: out<=0;
   2413: out<=0;
   2414: out<=0;
   2415: out<=0;
   2416: out<=0;
   2417: out<=1;
   2418: out<=0;
   2419: out<=1;
   2420: out<=1;
   2421: out<=1;
   2422: out<=0;
   2423: out<=0;
   2424: out<=0;
   2425: out<=0;
   2426: out<=0;
   2427: out<=0;
   2428: out<=1;
   2429: out<=0;
   2430: out<=0;
   2431: out<=1;
   2432: out<=1;
   2433: out<=0;
   2434: out<=0;
   2435: out<=1;
   2436: out<=0;
   2437: out<=0;
   2438: out<=0;
   2439: out<=0;
   2440: out<=0;
   2441: out<=0;
   2442: out<=1;
   2443: out<=1;
   2444: out<=1;
   2445: out<=0;
   2446: out<=1;
   2447: out<=0;
   2448: out<=0;
   2449: out<=0;
   2450: out<=0;
   2451: out<=0;
   2452: out<=0;
   2453: out<=1;
   2454: out<=1;
   2455: out<=0;
   2456: out<=0;
   2457: out<=1;
   2458: out<=0;
   2459: out<=1;
   2460: out<=0;
   2461: out<=0;
   2462: out<=1;
   2463: out<=1;
   2464: out<=0;
   2465: out<=0;
   2466: out<=1;
   2467: out<=1;
   2468: out<=0;
   2469: out<=1;
   2470: out<=0;
   2471: out<=1;
   2472: out<=1;
   2473: out<=0;
   2474: out<=0;
   2475: out<=1;
   2476: out<=1;
   2477: out<=1;
   2478: out<=1;
   2479: out<=1;
   2480: out<=1;
   2481: out<=0;
   2482: out<=1;
   2483: out<=0;
   2484: out<=0;
   2485: out<=0;
   2486: out<=1;
   2487: out<=1;
   2488: out<=1;
   2489: out<=1;
   2490: out<=1;
   2491: out<=1;
   2492: out<=0;
   2493: out<=1;
   2494: out<=1;
   2495: out<=0;
   2496: out<=0;
   2497: out<=1;
   2498: out<=1;
   2499: out<=0;
   2500: out<=1;
   2501: out<=1;
   2502: out<=1;
   2503: out<=1;
   2504: out<=1;
   2505: out<=1;
   2506: out<=0;
   2507: out<=0;
   2508: out<=0;
   2509: out<=1;
   2510: out<=0;
   2511: out<=1;
   2512: out<=0;
   2513: out<=0;
   2514: out<=0;
   2515: out<=0;
   2516: out<=0;
   2517: out<=1;
   2518: out<=1;
   2519: out<=0;
   2520: out<=0;
   2521: out<=1;
   2522: out<=0;
   2523: out<=1;
   2524: out<=0;
   2525: out<=0;
   2526: out<=1;
   2527: out<=1;
   2528: out<=0;
   2529: out<=0;
   2530: out<=1;
   2531: out<=1;
   2532: out<=0;
   2533: out<=1;
   2534: out<=0;
   2535: out<=1;
   2536: out<=1;
   2537: out<=0;
   2538: out<=0;
   2539: out<=1;
   2540: out<=1;
   2541: out<=1;
   2542: out<=1;
   2543: out<=1;
   2544: out<=0;
   2545: out<=1;
   2546: out<=0;
   2547: out<=1;
   2548: out<=1;
   2549: out<=1;
   2550: out<=0;
   2551: out<=0;
   2552: out<=0;
   2553: out<=0;
   2554: out<=0;
   2555: out<=0;
   2556: out<=1;
   2557: out<=0;
   2558: out<=0;
   2559: out<=1;
   2560: out<=0;
   2561: out<=1;
   2562: out<=0;
   2563: out<=1;
   2564: out<=1;
   2565: out<=1;
   2566: out<=0;
   2567: out<=0;
   2568: out<=0;
   2569: out<=0;
   2570: out<=0;
   2571: out<=0;
   2572: out<=1;
   2573: out<=0;
   2574: out<=0;
   2575: out<=1;
   2576: out<=0;
   2577: out<=0;
   2578: out<=1;
   2579: out<=1;
   2580: out<=0;
   2581: out<=1;
   2582: out<=0;
   2583: out<=1;
   2584: out<=1;
   2585: out<=0;
   2586: out<=0;
   2587: out<=1;
   2588: out<=1;
   2589: out<=1;
   2590: out<=1;
   2591: out<=1;
   2592: out<=0;
   2593: out<=0;
   2594: out<=0;
   2595: out<=0;
   2596: out<=0;
   2597: out<=1;
   2598: out<=1;
   2599: out<=0;
   2600: out<=0;
   2601: out<=1;
   2602: out<=0;
   2603: out<=1;
   2604: out<=0;
   2605: out<=0;
   2606: out<=1;
   2607: out<=1;
   2608: out<=0;
   2609: out<=1;
   2610: out<=1;
   2611: out<=0;
   2612: out<=1;
   2613: out<=1;
   2614: out<=1;
   2615: out<=1;
   2616: out<=1;
   2617: out<=1;
   2618: out<=0;
   2619: out<=0;
   2620: out<=0;
   2621: out<=1;
   2622: out<=0;
   2623: out<=1;
   2624: out<=1;
   2625: out<=0;
   2626: out<=1;
   2627: out<=0;
   2628: out<=0;
   2629: out<=0;
   2630: out<=1;
   2631: out<=1;
   2632: out<=1;
   2633: out<=1;
   2634: out<=1;
   2635: out<=1;
   2636: out<=0;
   2637: out<=1;
   2638: out<=1;
   2639: out<=0;
   2640: out<=0;
   2641: out<=0;
   2642: out<=1;
   2643: out<=1;
   2644: out<=0;
   2645: out<=1;
   2646: out<=0;
   2647: out<=1;
   2648: out<=1;
   2649: out<=0;
   2650: out<=0;
   2651: out<=1;
   2652: out<=1;
   2653: out<=1;
   2654: out<=1;
   2655: out<=1;
   2656: out<=0;
   2657: out<=0;
   2658: out<=0;
   2659: out<=0;
   2660: out<=0;
   2661: out<=1;
   2662: out<=1;
   2663: out<=0;
   2664: out<=0;
   2665: out<=1;
   2666: out<=0;
   2667: out<=1;
   2668: out<=0;
   2669: out<=0;
   2670: out<=1;
   2671: out<=1;
   2672: out<=1;
   2673: out<=0;
   2674: out<=0;
   2675: out<=1;
   2676: out<=0;
   2677: out<=0;
   2678: out<=0;
   2679: out<=0;
   2680: out<=0;
   2681: out<=0;
   2682: out<=1;
   2683: out<=1;
   2684: out<=1;
   2685: out<=0;
   2686: out<=1;
   2687: out<=0;
   2688: out<=0;
   2689: out<=1;
   2690: out<=0;
   2691: out<=1;
   2692: out<=1;
   2693: out<=1;
   2694: out<=0;
   2695: out<=0;
   2696: out<=0;
   2697: out<=0;
   2698: out<=0;
   2699: out<=0;
   2700: out<=1;
   2701: out<=0;
   2702: out<=0;
   2703: out<=1;
   2704: out<=1;
   2705: out<=1;
   2706: out<=0;
   2707: out<=0;
   2708: out<=1;
   2709: out<=0;
   2710: out<=1;
   2711: out<=0;
   2712: out<=0;
   2713: out<=1;
   2714: out<=1;
   2715: out<=0;
   2716: out<=0;
   2717: out<=0;
   2718: out<=0;
   2719: out<=0;
   2720: out<=0;
   2721: out<=0;
   2722: out<=0;
   2723: out<=0;
   2724: out<=0;
   2725: out<=1;
   2726: out<=1;
   2727: out<=0;
   2728: out<=0;
   2729: out<=1;
   2730: out<=0;
   2731: out<=1;
   2732: out<=0;
   2733: out<=0;
   2734: out<=1;
   2735: out<=1;
   2736: out<=1;
   2737: out<=0;
   2738: out<=0;
   2739: out<=1;
   2740: out<=0;
   2741: out<=0;
   2742: out<=0;
   2743: out<=0;
   2744: out<=0;
   2745: out<=0;
   2746: out<=1;
   2747: out<=1;
   2748: out<=1;
   2749: out<=0;
   2750: out<=1;
   2751: out<=0;
   2752: out<=1;
   2753: out<=0;
   2754: out<=1;
   2755: out<=0;
   2756: out<=0;
   2757: out<=0;
   2758: out<=1;
   2759: out<=1;
   2760: out<=1;
   2761: out<=1;
   2762: out<=1;
   2763: out<=1;
   2764: out<=0;
   2765: out<=1;
   2766: out<=1;
   2767: out<=0;
   2768: out<=1;
   2769: out<=1;
   2770: out<=0;
   2771: out<=0;
   2772: out<=1;
   2773: out<=0;
   2774: out<=1;
   2775: out<=0;
   2776: out<=0;
   2777: out<=1;
   2778: out<=1;
   2779: out<=0;
   2780: out<=0;
   2781: out<=0;
   2782: out<=0;
   2783: out<=0;
   2784: out<=0;
   2785: out<=0;
   2786: out<=0;
   2787: out<=0;
   2788: out<=0;
   2789: out<=1;
   2790: out<=1;
   2791: out<=0;
   2792: out<=0;
   2793: out<=1;
   2794: out<=0;
   2795: out<=1;
   2796: out<=0;
   2797: out<=0;
   2798: out<=1;
   2799: out<=1;
   2800: out<=0;
   2801: out<=1;
   2802: out<=1;
   2803: out<=0;
   2804: out<=1;
   2805: out<=1;
   2806: out<=1;
   2807: out<=1;
   2808: out<=1;
   2809: out<=1;
   2810: out<=0;
   2811: out<=0;
   2812: out<=0;
   2813: out<=1;
   2814: out<=0;
   2815: out<=1;
   2816: out<=0;
   2817: out<=0;
   2818: out<=1;
   2819: out<=1;
   2820: out<=0;
   2821: out<=1;
   2822: out<=0;
   2823: out<=1;
   2824: out<=1;
   2825: out<=0;
   2826: out<=0;
   2827: out<=1;
   2828: out<=1;
   2829: out<=1;
   2830: out<=1;
   2831: out<=1;
   2832: out<=1;
   2833: out<=0;
   2834: out<=1;
   2835: out<=0;
   2836: out<=0;
   2837: out<=0;
   2838: out<=1;
   2839: out<=1;
   2840: out<=1;
   2841: out<=1;
   2842: out<=1;
   2843: out<=1;
   2844: out<=0;
   2845: out<=1;
   2846: out<=1;
   2847: out<=0;
   2848: out<=1;
   2849: out<=0;
   2850: out<=0;
   2851: out<=1;
   2852: out<=0;
   2853: out<=0;
   2854: out<=0;
   2855: out<=0;
   2856: out<=0;
   2857: out<=0;
   2858: out<=1;
   2859: out<=1;
   2860: out<=1;
   2861: out<=0;
   2862: out<=1;
   2863: out<=0;
   2864: out<=0;
   2865: out<=0;
   2866: out<=0;
   2867: out<=0;
   2868: out<=0;
   2869: out<=1;
   2870: out<=1;
   2871: out<=0;
   2872: out<=0;
   2873: out<=1;
   2874: out<=0;
   2875: out<=1;
   2876: out<=0;
   2877: out<=0;
   2878: out<=1;
   2879: out<=1;
   2880: out<=0;
   2881: out<=0;
   2882: out<=1;
   2883: out<=1;
   2884: out<=0;
   2885: out<=1;
   2886: out<=0;
   2887: out<=1;
   2888: out<=1;
   2889: out<=0;
   2890: out<=0;
   2891: out<=1;
   2892: out<=1;
   2893: out<=1;
   2894: out<=1;
   2895: out<=1;
   2896: out<=0;
   2897: out<=1;
   2898: out<=0;
   2899: out<=1;
   2900: out<=1;
   2901: out<=1;
   2902: out<=0;
   2903: out<=0;
   2904: out<=0;
   2905: out<=0;
   2906: out<=0;
   2907: out<=0;
   2908: out<=1;
   2909: out<=0;
   2910: out<=0;
   2911: out<=1;
   2912: out<=0;
   2913: out<=1;
   2914: out<=1;
   2915: out<=0;
   2916: out<=1;
   2917: out<=1;
   2918: out<=1;
   2919: out<=1;
   2920: out<=1;
   2921: out<=1;
   2922: out<=0;
   2923: out<=0;
   2924: out<=0;
   2925: out<=1;
   2926: out<=0;
   2927: out<=1;
   2928: out<=0;
   2929: out<=0;
   2930: out<=0;
   2931: out<=0;
   2932: out<=0;
   2933: out<=1;
   2934: out<=1;
   2935: out<=0;
   2936: out<=0;
   2937: out<=1;
   2938: out<=0;
   2939: out<=1;
   2940: out<=0;
   2941: out<=0;
   2942: out<=1;
   2943: out<=1;
   2944: out<=1;
   2945: out<=1;
   2946: out<=0;
   2947: out<=0;
   2948: out<=1;
   2949: out<=0;
   2950: out<=1;
   2951: out<=0;
   2952: out<=0;
   2953: out<=1;
   2954: out<=1;
   2955: out<=0;
   2956: out<=0;
   2957: out<=0;
   2958: out<=0;
   2959: out<=0;
   2960: out<=1;
   2961: out<=0;
   2962: out<=1;
   2963: out<=0;
   2964: out<=0;
   2965: out<=0;
   2966: out<=1;
   2967: out<=1;
   2968: out<=1;
   2969: out<=1;
   2970: out<=1;
   2971: out<=1;
   2972: out<=0;
   2973: out<=1;
   2974: out<=1;
   2975: out<=0;
   2976: out<=0;
   2977: out<=1;
   2978: out<=1;
   2979: out<=0;
   2980: out<=1;
   2981: out<=1;
   2982: out<=1;
   2983: out<=1;
   2984: out<=1;
   2985: out<=1;
   2986: out<=0;
   2987: out<=0;
   2988: out<=0;
   2989: out<=1;
   2990: out<=0;
   2991: out<=1;
   2992: out<=0;
   2993: out<=0;
   2994: out<=0;
   2995: out<=0;
   2996: out<=0;
   2997: out<=1;
   2998: out<=1;
   2999: out<=0;
   3000: out<=0;
   3001: out<=1;
   3002: out<=0;
   3003: out<=1;
   3004: out<=0;
   3005: out<=0;
   3006: out<=1;
   3007: out<=1;
   3008: out<=1;
   3009: out<=1;
   3010: out<=0;
   3011: out<=0;
   3012: out<=1;
   3013: out<=0;
   3014: out<=1;
   3015: out<=0;
   3016: out<=0;
   3017: out<=1;
   3018: out<=1;
   3019: out<=0;
   3020: out<=0;
   3021: out<=0;
   3022: out<=0;
   3023: out<=0;
   3024: out<=0;
   3025: out<=1;
   3026: out<=0;
   3027: out<=1;
   3028: out<=1;
   3029: out<=1;
   3030: out<=0;
   3031: out<=0;
   3032: out<=0;
   3033: out<=0;
   3034: out<=0;
   3035: out<=0;
   3036: out<=1;
   3037: out<=0;
   3038: out<=0;
   3039: out<=1;
   3040: out<=1;
   3041: out<=0;
   3042: out<=0;
   3043: out<=1;
   3044: out<=0;
   3045: out<=0;
   3046: out<=0;
   3047: out<=0;
   3048: out<=0;
   3049: out<=0;
   3050: out<=1;
   3051: out<=1;
   3052: out<=1;
   3053: out<=0;
   3054: out<=1;
   3055: out<=0;
   3056: out<=0;
   3057: out<=0;
   3058: out<=0;
   3059: out<=0;
   3060: out<=0;
   3061: out<=1;
   3062: out<=1;
   3063: out<=0;
   3064: out<=0;
   3065: out<=1;
   3066: out<=0;
   3067: out<=1;
   3068: out<=0;
   3069: out<=0;
   3070: out<=1;
   3071: out<=1;
   3072: out<=1;
   3073: out<=0;
   3074: out<=0;
   3075: out<=1;
   3076: out<=1;
   3077: out<=1;
   3078: out<=1;
   3079: out<=1;
   3080: out<=1;
   3081: out<=1;
   3082: out<=0;
   3083: out<=0;
   3084: out<=1;
   3085: out<=0;
   3086: out<=1;
   3087: out<=0;
   3088: out<=0;
   3089: out<=0;
   3090: out<=0;
   3091: out<=0;
   3092: out<=1;
   3093: out<=0;
   3094: out<=0;
   3095: out<=1;
   3096: out<=1;
   3097: out<=0;
   3098: out<=1;
   3099: out<=0;
   3100: out<=0;
   3101: out<=0;
   3102: out<=1;
   3103: out<=1;
   3104: out<=1;
   3105: out<=1;
   3106: out<=0;
   3107: out<=0;
   3108: out<=0;
   3109: out<=1;
   3110: out<=0;
   3111: out<=1;
   3112: out<=1;
   3113: out<=0;
   3114: out<=0;
   3115: out<=1;
   3116: out<=0;
   3117: out<=0;
   3118: out<=0;
   3119: out<=0;
   3120: out<=0;
   3121: out<=1;
   3122: out<=0;
   3123: out<=1;
   3124: out<=0;
   3125: out<=0;
   3126: out<=1;
   3127: out<=1;
   3128: out<=1;
   3129: out<=1;
   3130: out<=1;
   3131: out<=1;
   3132: out<=1;
   3133: out<=0;
   3134: out<=0;
   3135: out<=1;
   3136: out<=0;
   3137: out<=1;
   3138: out<=1;
   3139: out<=0;
   3140: out<=0;
   3141: out<=0;
   3142: out<=0;
   3143: out<=0;
   3144: out<=0;
   3145: out<=0;
   3146: out<=1;
   3147: out<=1;
   3148: out<=0;
   3149: out<=1;
   3150: out<=0;
   3151: out<=1;
   3152: out<=0;
   3153: out<=0;
   3154: out<=0;
   3155: out<=0;
   3156: out<=1;
   3157: out<=0;
   3158: out<=0;
   3159: out<=1;
   3160: out<=1;
   3161: out<=0;
   3162: out<=1;
   3163: out<=0;
   3164: out<=0;
   3165: out<=0;
   3166: out<=1;
   3167: out<=1;
   3168: out<=1;
   3169: out<=1;
   3170: out<=0;
   3171: out<=0;
   3172: out<=0;
   3173: out<=1;
   3174: out<=0;
   3175: out<=1;
   3176: out<=1;
   3177: out<=0;
   3178: out<=0;
   3179: out<=1;
   3180: out<=0;
   3181: out<=0;
   3182: out<=0;
   3183: out<=0;
   3184: out<=1;
   3185: out<=0;
   3186: out<=1;
   3187: out<=0;
   3188: out<=1;
   3189: out<=1;
   3190: out<=0;
   3191: out<=0;
   3192: out<=0;
   3193: out<=0;
   3194: out<=0;
   3195: out<=0;
   3196: out<=0;
   3197: out<=1;
   3198: out<=1;
   3199: out<=0;
   3200: out<=0;
   3201: out<=1;
   3202: out<=1;
   3203: out<=0;
   3204: out<=0;
   3205: out<=0;
   3206: out<=0;
   3207: out<=0;
   3208: out<=0;
   3209: out<=0;
   3210: out<=1;
   3211: out<=1;
   3212: out<=0;
   3213: out<=1;
   3214: out<=0;
   3215: out<=1;
   3216: out<=0;
   3217: out<=0;
   3218: out<=0;
   3219: out<=0;
   3220: out<=1;
   3221: out<=0;
   3222: out<=0;
   3223: out<=1;
   3224: out<=1;
   3225: out<=0;
   3226: out<=1;
   3227: out<=0;
   3228: out<=0;
   3229: out<=0;
   3230: out<=1;
   3231: out<=1;
   3232: out<=0;
   3233: out<=0;
   3234: out<=1;
   3235: out<=1;
   3236: out<=1;
   3237: out<=0;
   3238: out<=1;
   3239: out<=0;
   3240: out<=0;
   3241: out<=1;
   3242: out<=1;
   3243: out<=0;
   3244: out<=1;
   3245: out<=1;
   3246: out<=1;
   3247: out<=1;
   3248: out<=0;
   3249: out<=1;
   3250: out<=0;
   3251: out<=1;
   3252: out<=0;
   3253: out<=0;
   3254: out<=1;
   3255: out<=1;
   3256: out<=1;
   3257: out<=1;
   3258: out<=1;
   3259: out<=1;
   3260: out<=1;
   3261: out<=0;
   3262: out<=0;
   3263: out<=1;
   3264: out<=1;
   3265: out<=0;
   3266: out<=0;
   3267: out<=1;
   3268: out<=1;
   3269: out<=1;
   3270: out<=1;
   3271: out<=1;
   3272: out<=1;
   3273: out<=1;
   3274: out<=0;
   3275: out<=0;
   3276: out<=1;
   3277: out<=0;
   3278: out<=1;
   3279: out<=0;
   3280: out<=0;
   3281: out<=0;
   3282: out<=0;
   3283: out<=0;
   3284: out<=1;
   3285: out<=0;
   3286: out<=0;
   3287: out<=1;
   3288: out<=1;
   3289: out<=0;
   3290: out<=1;
   3291: out<=0;
   3292: out<=0;
   3293: out<=0;
   3294: out<=1;
   3295: out<=1;
   3296: out<=0;
   3297: out<=0;
   3298: out<=1;
   3299: out<=1;
   3300: out<=1;
   3301: out<=0;
   3302: out<=1;
   3303: out<=0;
   3304: out<=0;
   3305: out<=1;
   3306: out<=1;
   3307: out<=0;
   3308: out<=1;
   3309: out<=1;
   3310: out<=1;
   3311: out<=1;
   3312: out<=1;
   3313: out<=0;
   3314: out<=1;
   3315: out<=0;
   3316: out<=1;
   3317: out<=1;
   3318: out<=0;
   3319: out<=0;
   3320: out<=0;
   3321: out<=0;
   3322: out<=0;
   3323: out<=0;
   3324: out<=0;
   3325: out<=1;
   3326: out<=1;
   3327: out<=0;
   3328: out<=0;
   3329: out<=0;
   3330: out<=0;
   3331: out<=0;
   3332: out<=1;
   3333: out<=0;
   3334: out<=0;
   3335: out<=1;
   3336: out<=1;
   3337: out<=0;
   3338: out<=1;
   3339: out<=0;
   3340: out<=0;
   3341: out<=0;
   3342: out<=1;
   3343: out<=1;
   3344: out<=0;
   3345: out<=1;
   3346: out<=1;
   3347: out<=0;
   3348: out<=0;
   3349: out<=0;
   3350: out<=0;
   3351: out<=0;
   3352: out<=0;
   3353: out<=0;
   3354: out<=1;
   3355: out<=1;
   3356: out<=0;
   3357: out<=1;
   3358: out<=0;
   3359: out<=1;
   3360: out<=1;
   3361: out<=0;
   3362: out<=1;
   3363: out<=0;
   3364: out<=1;
   3365: out<=1;
   3366: out<=0;
   3367: out<=0;
   3368: out<=0;
   3369: out<=0;
   3370: out<=0;
   3371: out<=0;
   3372: out<=0;
   3373: out<=1;
   3374: out<=1;
   3375: out<=0;
   3376: out<=1;
   3377: out<=1;
   3378: out<=0;
   3379: out<=0;
   3380: out<=0;
   3381: out<=1;
   3382: out<=0;
   3383: out<=1;
   3384: out<=1;
   3385: out<=0;
   3386: out<=0;
   3387: out<=1;
   3388: out<=0;
   3389: out<=0;
   3390: out<=0;
   3391: out<=0;
   3392: out<=0;
   3393: out<=0;
   3394: out<=0;
   3395: out<=0;
   3396: out<=1;
   3397: out<=0;
   3398: out<=0;
   3399: out<=1;
   3400: out<=1;
   3401: out<=0;
   3402: out<=1;
   3403: out<=0;
   3404: out<=0;
   3405: out<=0;
   3406: out<=1;
   3407: out<=1;
   3408: out<=1;
   3409: out<=0;
   3410: out<=0;
   3411: out<=1;
   3412: out<=1;
   3413: out<=1;
   3414: out<=1;
   3415: out<=1;
   3416: out<=1;
   3417: out<=1;
   3418: out<=0;
   3419: out<=0;
   3420: out<=1;
   3421: out<=0;
   3422: out<=1;
   3423: out<=0;
   3424: out<=0;
   3425: out<=1;
   3426: out<=0;
   3427: out<=1;
   3428: out<=0;
   3429: out<=0;
   3430: out<=1;
   3431: out<=1;
   3432: out<=1;
   3433: out<=1;
   3434: out<=1;
   3435: out<=1;
   3436: out<=1;
   3437: out<=0;
   3438: out<=0;
   3439: out<=1;
   3440: out<=1;
   3441: out<=1;
   3442: out<=0;
   3443: out<=0;
   3444: out<=0;
   3445: out<=1;
   3446: out<=0;
   3447: out<=1;
   3448: out<=1;
   3449: out<=0;
   3450: out<=0;
   3451: out<=1;
   3452: out<=0;
   3453: out<=0;
   3454: out<=0;
   3455: out<=0;
   3456: out<=0;
   3457: out<=0;
   3458: out<=0;
   3459: out<=0;
   3460: out<=1;
   3461: out<=0;
   3462: out<=0;
   3463: out<=1;
   3464: out<=1;
   3465: out<=0;
   3466: out<=1;
   3467: out<=0;
   3468: out<=0;
   3469: out<=0;
   3470: out<=1;
   3471: out<=1;
   3472: out<=1;
   3473: out<=0;
   3474: out<=0;
   3475: out<=1;
   3476: out<=1;
   3477: out<=1;
   3478: out<=1;
   3479: out<=1;
   3480: out<=1;
   3481: out<=1;
   3482: out<=0;
   3483: out<=0;
   3484: out<=1;
   3485: out<=0;
   3486: out<=1;
   3487: out<=0;
   3488: out<=1;
   3489: out<=0;
   3490: out<=1;
   3491: out<=0;
   3492: out<=1;
   3493: out<=1;
   3494: out<=0;
   3495: out<=0;
   3496: out<=0;
   3497: out<=0;
   3498: out<=0;
   3499: out<=0;
   3500: out<=0;
   3501: out<=1;
   3502: out<=1;
   3503: out<=0;
   3504: out<=0;
   3505: out<=0;
   3506: out<=1;
   3507: out<=1;
   3508: out<=1;
   3509: out<=0;
   3510: out<=1;
   3511: out<=0;
   3512: out<=0;
   3513: out<=1;
   3514: out<=1;
   3515: out<=0;
   3516: out<=1;
   3517: out<=1;
   3518: out<=1;
   3519: out<=1;
   3520: out<=0;
   3521: out<=0;
   3522: out<=0;
   3523: out<=0;
   3524: out<=1;
   3525: out<=0;
   3526: out<=0;
   3527: out<=1;
   3528: out<=1;
   3529: out<=0;
   3530: out<=1;
   3531: out<=0;
   3532: out<=0;
   3533: out<=0;
   3534: out<=1;
   3535: out<=1;
   3536: out<=0;
   3537: out<=1;
   3538: out<=1;
   3539: out<=0;
   3540: out<=0;
   3541: out<=0;
   3542: out<=0;
   3543: out<=0;
   3544: out<=0;
   3545: out<=0;
   3546: out<=1;
   3547: out<=1;
   3548: out<=0;
   3549: out<=1;
   3550: out<=0;
   3551: out<=1;
   3552: out<=0;
   3553: out<=1;
   3554: out<=0;
   3555: out<=1;
   3556: out<=0;
   3557: out<=0;
   3558: out<=1;
   3559: out<=1;
   3560: out<=1;
   3561: out<=1;
   3562: out<=1;
   3563: out<=1;
   3564: out<=1;
   3565: out<=0;
   3566: out<=0;
   3567: out<=1;
   3568: out<=0;
   3569: out<=0;
   3570: out<=1;
   3571: out<=1;
   3572: out<=1;
   3573: out<=0;
   3574: out<=1;
   3575: out<=0;
   3576: out<=0;
   3577: out<=1;
   3578: out<=1;
   3579: out<=0;
   3580: out<=1;
   3581: out<=1;
   3582: out<=1;
   3583: out<=1;
   3584: out<=0;
   3585: out<=0;
   3586: out<=1;
   3587: out<=1;
   3588: out<=1;
   3589: out<=0;
   3590: out<=1;
   3591: out<=0;
   3592: out<=0;
   3593: out<=1;
   3594: out<=1;
   3595: out<=0;
   3596: out<=1;
   3597: out<=1;
   3598: out<=1;
   3599: out<=1;
   3600: out<=0;
   3601: out<=1;
   3602: out<=0;
   3603: out<=1;
   3604: out<=0;
   3605: out<=0;
   3606: out<=1;
   3607: out<=1;
   3608: out<=1;
   3609: out<=1;
   3610: out<=1;
   3611: out<=1;
   3612: out<=1;
   3613: out<=0;
   3614: out<=0;
   3615: out<=1;
   3616: out<=0;
   3617: out<=1;
   3618: out<=1;
   3619: out<=0;
   3620: out<=0;
   3621: out<=0;
   3622: out<=0;
   3623: out<=0;
   3624: out<=0;
   3625: out<=0;
   3626: out<=1;
   3627: out<=1;
   3628: out<=0;
   3629: out<=1;
   3630: out<=0;
   3631: out<=1;
   3632: out<=0;
   3633: out<=0;
   3634: out<=0;
   3635: out<=0;
   3636: out<=1;
   3637: out<=0;
   3638: out<=0;
   3639: out<=1;
   3640: out<=1;
   3641: out<=0;
   3642: out<=1;
   3643: out<=0;
   3644: out<=0;
   3645: out<=0;
   3646: out<=1;
   3647: out<=1;
   3648: out<=0;
   3649: out<=0;
   3650: out<=1;
   3651: out<=1;
   3652: out<=1;
   3653: out<=0;
   3654: out<=1;
   3655: out<=0;
   3656: out<=0;
   3657: out<=1;
   3658: out<=1;
   3659: out<=0;
   3660: out<=1;
   3661: out<=1;
   3662: out<=1;
   3663: out<=1;
   3664: out<=1;
   3665: out<=0;
   3666: out<=1;
   3667: out<=0;
   3668: out<=1;
   3669: out<=1;
   3670: out<=0;
   3671: out<=0;
   3672: out<=0;
   3673: out<=0;
   3674: out<=0;
   3675: out<=0;
   3676: out<=0;
   3677: out<=1;
   3678: out<=1;
   3679: out<=0;
   3680: out<=1;
   3681: out<=0;
   3682: out<=0;
   3683: out<=1;
   3684: out<=1;
   3685: out<=1;
   3686: out<=1;
   3687: out<=1;
   3688: out<=1;
   3689: out<=1;
   3690: out<=0;
   3691: out<=0;
   3692: out<=1;
   3693: out<=0;
   3694: out<=1;
   3695: out<=0;
   3696: out<=0;
   3697: out<=0;
   3698: out<=0;
   3699: out<=0;
   3700: out<=1;
   3701: out<=0;
   3702: out<=0;
   3703: out<=1;
   3704: out<=1;
   3705: out<=0;
   3706: out<=1;
   3707: out<=0;
   3708: out<=0;
   3709: out<=0;
   3710: out<=1;
   3711: out<=1;
   3712: out<=1;
   3713: out<=1;
   3714: out<=0;
   3715: out<=0;
   3716: out<=0;
   3717: out<=1;
   3718: out<=0;
   3719: out<=1;
   3720: out<=1;
   3721: out<=0;
   3722: out<=0;
   3723: out<=1;
   3724: out<=0;
   3725: out<=0;
   3726: out<=0;
   3727: out<=0;
   3728: out<=0;
   3729: out<=1;
   3730: out<=0;
   3731: out<=1;
   3732: out<=0;
   3733: out<=0;
   3734: out<=1;
   3735: out<=1;
   3736: out<=1;
   3737: out<=1;
   3738: out<=1;
   3739: out<=1;
   3740: out<=1;
   3741: out<=0;
   3742: out<=0;
   3743: out<=1;
   3744: out<=1;
   3745: out<=0;
   3746: out<=0;
   3747: out<=1;
   3748: out<=1;
   3749: out<=1;
   3750: out<=1;
   3751: out<=1;
   3752: out<=1;
   3753: out<=1;
   3754: out<=0;
   3755: out<=0;
   3756: out<=1;
   3757: out<=0;
   3758: out<=1;
   3759: out<=0;
   3760: out<=0;
   3761: out<=0;
   3762: out<=0;
   3763: out<=0;
   3764: out<=1;
   3765: out<=0;
   3766: out<=0;
   3767: out<=1;
   3768: out<=1;
   3769: out<=0;
   3770: out<=1;
   3771: out<=0;
   3772: out<=0;
   3773: out<=0;
   3774: out<=1;
   3775: out<=1;
   3776: out<=1;
   3777: out<=1;
   3778: out<=0;
   3779: out<=0;
   3780: out<=0;
   3781: out<=1;
   3782: out<=0;
   3783: out<=1;
   3784: out<=1;
   3785: out<=0;
   3786: out<=0;
   3787: out<=1;
   3788: out<=0;
   3789: out<=0;
   3790: out<=0;
   3791: out<=0;
   3792: out<=1;
   3793: out<=0;
   3794: out<=1;
   3795: out<=0;
   3796: out<=1;
   3797: out<=1;
   3798: out<=0;
   3799: out<=0;
   3800: out<=0;
   3801: out<=0;
   3802: out<=0;
   3803: out<=0;
   3804: out<=0;
   3805: out<=1;
   3806: out<=1;
   3807: out<=0;
   3808: out<=0;
   3809: out<=1;
   3810: out<=1;
   3811: out<=0;
   3812: out<=0;
   3813: out<=0;
   3814: out<=0;
   3815: out<=0;
   3816: out<=0;
   3817: out<=0;
   3818: out<=1;
   3819: out<=1;
   3820: out<=0;
   3821: out<=1;
   3822: out<=0;
   3823: out<=1;
   3824: out<=0;
   3825: out<=0;
   3826: out<=0;
   3827: out<=0;
   3828: out<=1;
   3829: out<=0;
   3830: out<=0;
   3831: out<=1;
   3832: out<=1;
   3833: out<=0;
   3834: out<=1;
   3835: out<=0;
   3836: out<=0;
   3837: out<=0;
   3838: out<=1;
   3839: out<=1;
   3840: out<=1;
   3841: out<=0;
   3842: out<=1;
   3843: out<=0;
   3844: out<=1;
   3845: out<=1;
   3846: out<=0;
   3847: out<=0;
   3848: out<=0;
   3849: out<=0;
   3850: out<=0;
   3851: out<=0;
   3852: out<=0;
   3853: out<=1;
   3854: out<=1;
   3855: out<=0;
   3856: out<=0;
   3857: out<=0;
   3858: out<=1;
   3859: out<=1;
   3860: out<=1;
   3861: out<=0;
   3862: out<=1;
   3863: out<=0;
   3864: out<=0;
   3865: out<=1;
   3866: out<=1;
   3867: out<=0;
   3868: out<=1;
   3869: out<=1;
   3870: out<=1;
   3871: out<=1;
   3872: out<=0;
   3873: out<=0;
   3874: out<=0;
   3875: out<=0;
   3876: out<=1;
   3877: out<=0;
   3878: out<=0;
   3879: out<=1;
   3880: out<=1;
   3881: out<=0;
   3882: out<=1;
   3883: out<=0;
   3884: out<=0;
   3885: out<=0;
   3886: out<=1;
   3887: out<=1;
   3888: out<=1;
   3889: out<=0;
   3890: out<=0;
   3891: out<=1;
   3892: out<=1;
   3893: out<=1;
   3894: out<=1;
   3895: out<=1;
   3896: out<=1;
   3897: out<=1;
   3898: out<=0;
   3899: out<=0;
   3900: out<=1;
   3901: out<=0;
   3902: out<=1;
   3903: out<=0;
   3904: out<=0;
   3905: out<=1;
   3906: out<=0;
   3907: out<=1;
   3908: out<=0;
   3909: out<=0;
   3910: out<=1;
   3911: out<=1;
   3912: out<=1;
   3913: out<=1;
   3914: out<=1;
   3915: out<=1;
   3916: out<=1;
   3917: out<=0;
   3918: out<=0;
   3919: out<=1;
   3920: out<=0;
   3921: out<=0;
   3922: out<=1;
   3923: out<=1;
   3924: out<=1;
   3925: out<=0;
   3926: out<=1;
   3927: out<=0;
   3928: out<=0;
   3929: out<=1;
   3930: out<=1;
   3931: out<=0;
   3932: out<=1;
   3933: out<=1;
   3934: out<=1;
   3935: out<=1;
   3936: out<=0;
   3937: out<=0;
   3938: out<=0;
   3939: out<=0;
   3940: out<=1;
   3941: out<=0;
   3942: out<=0;
   3943: out<=1;
   3944: out<=1;
   3945: out<=0;
   3946: out<=1;
   3947: out<=0;
   3948: out<=0;
   3949: out<=0;
   3950: out<=1;
   3951: out<=1;
   3952: out<=0;
   3953: out<=1;
   3954: out<=1;
   3955: out<=0;
   3956: out<=0;
   3957: out<=0;
   3958: out<=0;
   3959: out<=0;
   3960: out<=0;
   3961: out<=0;
   3962: out<=1;
   3963: out<=1;
   3964: out<=0;
   3965: out<=1;
   3966: out<=0;
   3967: out<=1;
   3968: out<=1;
   3969: out<=0;
   3970: out<=1;
   3971: out<=0;
   3972: out<=1;
   3973: out<=1;
   3974: out<=0;
   3975: out<=0;
   3976: out<=0;
   3977: out<=0;
   3978: out<=0;
   3979: out<=0;
   3980: out<=0;
   3981: out<=1;
   3982: out<=1;
   3983: out<=0;
   3984: out<=1;
   3985: out<=1;
   3986: out<=0;
   3987: out<=0;
   3988: out<=0;
   3989: out<=1;
   3990: out<=0;
   3991: out<=1;
   3992: out<=1;
   3993: out<=0;
   3994: out<=0;
   3995: out<=1;
   3996: out<=0;
   3997: out<=0;
   3998: out<=0;
   3999: out<=0;
   4000: out<=0;
   4001: out<=0;
   4002: out<=0;
   4003: out<=0;
   4004: out<=1;
   4005: out<=0;
   4006: out<=0;
   4007: out<=1;
   4008: out<=1;
   4009: out<=0;
   4010: out<=1;
   4011: out<=0;
   4012: out<=0;
   4013: out<=0;
   4014: out<=1;
   4015: out<=1;
   4016: out<=0;
   4017: out<=1;
   4018: out<=1;
   4019: out<=0;
   4020: out<=0;
   4021: out<=0;
   4022: out<=0;
   4023: out<=0;
   4024: out<=0;
   4025: out<=0;
   4026: out<=1;
   4027: out<=1;
   4028: out<=0;
   4029: out<=1;
   4030: out<=0;
   4031: out<=1;
   4032: out<=0;
   4033: out<=1;
   4034: out<=0;
   4035: out<=1;
   4036: out<=0;
   4037: out<=0;
   4038: out<=1;
   4039: out<=1;
   4040: out<=1;
   4041: out<=1;
   4042: out<=1;
   4043: out<=1;
   4044: out<=1;
   4045: out<=0;
   4046: out<=0;
   4047: out<=1;
   4048: out<=1;
   4049: out<=1;
   4050: out<=0;
   4051: out<=0;
   4052: out<=0;
   4053: out<=1;
   4054: out<=0;
   4055: out<=1;
   4056: out<=1;
   4057: out<=0;
   4058: out<=0;
   4059: out<=1;
   4060: out<=0;
   4061: out<=0;
   4062: out<=0;
   4063: out<=0;
   4064: out<=0;
   4065: out<=0;
   4066: out<=0;
   4067: out<=0;
   4068: out<=1;
   4069: out<=0;
   4070: out<=0;
   4071: out<=1;
   4072: out<=1;
   4073: out<=0;
   4074: out<=1;
   4075: out<=0;
   4076: out<=0;
   4077: out<=0;
   4078: out<=1;
   4079: out<=1;
   4080: out<=1;
   4081: out<=0;
   4082: out<=0;
   4083: out<=1;
   4084: out<=1;
   4085: out<=1;
   4086: out<=1;
   4087: out<=1;
   4088: out<=1;
   4089: out<=1;
   4090: out<=0;
   4091: out<=0;
   4092: out<=1;
   4093: out<=0;
   4094: out<=1;
   4095: out<=0;
   4096: out<=1;
   4097: out<=0;
   4098: out<=1;
   4099: out<=0;
   4100: out<=0;
   4101: out<=0;
   4102: out<=1;
   4103: out<=1;
   4104: out<=0;
   4105: out<=0;
   4106: out<=0;
   4107: out<=0;
   4108: out<=1;
   4109: out<=0;
   4110: out<=0;
   4111: out<=1;
   4112: out<=0;
   4113: out<=0;
   4114: out<=1;
   4115: out<=1;
   4116: out<=0;
   4117: out<=1;
   4118: out<=0;
   4119: out<=1;
   4120: out<=0;
   4121: out<=1;
   4122: out<=1;
   4123: out<=0;
   4124: out<=0;
   4125: out<=0;
   4126: out<=0;
   4127: out<=0;
   4128: out<=1;
   4129: out<=1;
   4130: out<=1;
   4131: out<=1;
   4132: out<=1;
   4133: out<=0;
   4134: out<=0;
   4135: out<=1;
   4136: out<=0;
   4137: out<=1;
   4138: out<=0;
   4139: out<=1;
   4140: out<=0;
   4141: out<=0;
   4142: out<=1;
   4143: out<=1;
   4144: out<=0;
   4145: out<=1;
   4146: out<=1;
   4147: out<=0;
   4148: out<=1;
   4149: out<=1;
   4150: out<=1;
   4151: out<=1;
   4152: out<=0;
   4153: out<=0;
   4154: out<=1;
   4155: out<=1;
   4156: out<=1;
   4157: out<=0;
   4158: out<=1;
   4159: out<=0;
   4160: out<=0;
   4161: out<=1;
   4162: out<=0;
   4163: out<=1;
   4164: out<=1;
   4165: out<=1;
   4166: out<=0;
   4167: out<=0;
   4168: out<=1;
   4169: out<=1;
   4170: out<=1;
   4171: out<=1;
   4172: out<=0;
   4173: out<=1;
   4174: out<=1;
   4175: out<=0;
   4176: out<=0;
   4177: out<=0;
   4178: out<=1;
   4179: out<=1;
   4180: out<=0;
   4181: out<=1;
   4182: out<=0;
   4183: out<=1;
   4184: out<=0;
   4185: out<=1;
   4186: out<=1;
   4187: out<=0;
   4188: out<=0;
   4189: out<=0;
   4190: out<=0;
   4191: out<=0;
   4192: out<=1;
   4193: out<=1;
   4194: out<=1;
   4195: out<=1;
   4196: out<=1;
   4197: out<=0;
   4198: out<=0;
   4199: out<=1;
   4200: out<=0;
   4201: out<=1;
   4202: out<=0;
   4203: out<=1;
   4204: out<=0;
   4205: out<=0;
   4206: out<=1;
   4207: out<=1;
   4208: out<=1;
   4209: out<=0;
   4210: out<=0;
   4211: out<=1;
   4212: out<=0;
   4213: out<=0;
   4214: out<=0;
   4215: out<=0;
   4216: out<=1;
   4217: out<=1;
   4218: out<=0;
   4219: out<=0;
   4220: out<=0;
   4221: out<=1;
   4222: out<=0;
   4223: out<=1;
   4224: out<=1;
   4225: out<=0;
   4226: out<=1;
   4227: out<=0;
   4228: out<=0;
   4229: out<=0;
   4230: out<=1;
   4231: out<=1;
   4232: out<=0;
   4233: out<=0;
   4234: out<=0;
   4235: out<=0;
   4236: out<=1;
   4237: out<=0;
   4238: out<=0;
   4239: out<=1;
   4240: out<=1;
   4241: out<=1;
   4242: out<=0;
   4243: out<=0;
   4244: out<=1;
   4245: out<=0;
   4246: out<=1;
   4247: out<=0;
   4248: out<=1;
   4249: out<=0;
   4250: out<=0;
   4251: out<=1;
   4252: out<=1;
   4253: out<=1;
   4254: out<=1;
   4255: out<=1;
   4256: out<=1;
   4257: out<=1;
   4258: out<=1;
   4259: out<=1;
   4260: out<=1;
   4261: out<=0;
   4262: out<=0;
   4263: out<=1;
   4264: out<=0;
   4265: out<=1;
   4266: out<=0;
   4267: out<=1;
   4268: out<=0;
   4269: out<=0;
   4270: out<=1;
   4271: out<=1;
   4272: out<=1;
   4273: out<=0;
   4274: out<=0;
   4275: out<=1;
   4276: out<=0;
   4277: out<=0;
   4278: out<=0;
   4279: out<=0;
   4280: out<=1;
   4281: out<=1;
   4282: out<=0;
   4283: out<=0;
   4284: out<=0;
   4285: out<=1;
   4286: out<=0;
   4287: out<=1;
   4288: out<=0;
   4289: out<=1;
   4290: out<=0;
   4291: out<=1;
   4292: out<=1;
   4293: out<=1;
   4294: out<=0;
   4295: out<=0;
   4296: out<=1;
   4297: out<=1;
   4298: out<=1;
   4299: out<=1;
   4300: out<=0;
   4301: out<=1;
   4302: out<=1;
   4303: out<=0;
   4304: out<=1;
   4305: out<=1;
   4306: out<=0;
   4307: out<=0;
   4308: out<=1;
   4309: out<=0;
   4310: out<=1;
   4311: out<=0;
   4312: out<=1;
   4313: out<=0;
   4314: out<=0;
   4315: out<=1;
   4316: out<=1;
   4317: out<=1;
   4318: out<=1;
   4319: out<=1;
   4320: out<=1;
   4321: out<=1;
   4322: out<=1;
   4323: out<=1;
   4324: out<=1;
   4325: out<=0;
   4326: out<=0;
   4327: out<=1;
   4328: out<=0;
   4329: out<=1;
   4330: out<=0;
   4331: out<=1;
   4332: out<=0;
   4333: out<=0;
   4334: out<=1;
   4335: out<=1;
   4336: out<=0;
   4337: out<=1;
   4338: out<=1;
   4339: out<=0;
   4340: out<=1;
   4341: out<=1;
   4342: out<=1;
   4343: out<=1;
   4344: out<=0;
   4345: out<=0;
   4346: out<=1;
   4347: out<=1;
   4348: out<=1;
   4349: out<=0;
   4350: out<=1;
   4351: out<=0;
   4352: out<=0;
   4353: out<=0;
   4354: out<=1;
   4355: out<=1;
   4356: out<=0;
   4357: out<=1;
   4358: out<=0;
   4359: out<=1;
   4360: out<=0;
   4361: out<=1;
   4362: out<=1;
   4363: out<=0;
   4364: out<=0;
   4365: out<=0;
   4366: out<=0;
   4367: out<=0;
   4368: out<=0;
   4369: out<=1;
   4370: out<=0;
   4371: out<=1;
   4372: out<=1;
   4373: out<=1;
   4374: out<=0;
   4375: out<=0;
   4376: out<=1;
   4377: out<=1;
   4378: out<=1;
   4379: out<=1;
   4380: out<=0;
   4381: out<=1;
   4382: out<=1;
   4383: out<=0;
   4384: out<=1;
   4385: out<=0;
   4386: out<=0;
   4387: out<=1;
   4388: out<=0;
   4389: out<=0;
   4390: out<=0;
   4391: out<=0;
   4392: out<=1;
   4393: out<=1;
   4394: out<=0;
   4395: out<=0;
   4396: out<=0;
   4397: out<=1;
   4398: out<=0;
   4399: out<=1;
   4400: out<=1;
   4401: out<=1;
   4402: out<=1;
   4403: out<=1;
   4404: out<=1;
   4405: out<=0;
   4406: out<=0;
   4407: out<=1;
   4408: out<=0;
   4409: out<=1;
   4410: out<=0;
   4411: out<=1;
   4412: out<=0;
   4413: out<=0;
   4414: out<=1;
   4415: out<=1;
   4416: out<=0;
   4417: out<=0;
   4418: out<=1;
   4419: out<=1;
   4420: out<=0;
   4421: out<=1;
   4422: out<=0;
   4423: out<=1;
   4424: out<=0;
   4425: out<=1;
   4426: out<=1;
   4427: out<=0;
   4428: out<=0;
   4429: out<=0;
   4430: out<=0;
   4431: out<=0;
   4432: out<=1;
   4433: out<=0;
   4434: out<=1;
   4435: out<=0;
   4436: out<=0;
   4437: out<=0;
   4438: out<=1;
   4439: out<=1;
   4440: out<=0;
   4441: out<=0;
   4442: out<=0;
   4443: out<=0;
   4444: out<=1;
   4445: out<=0;
   4446: out<=0;
   4447: out<=1;
   4448: out<=0;
   4449: out<=1;
   4450: out<=1;
   4451: out<=0;
   4452: out<=1;
   4453: out<=1;
   4454: out<=1;
   4455: out<=1;
   4456: out<=0;
   4457: out<=0;
   4458: out<=1;
   4459: out<=1;
   4460: out<=1;
   4461: out<=0;
   4462: out<=1;
   4463: out<=0;
   4464: out<=1;
   4465: out<=1;
   4466: out<=1;
   4467: out<=1;
   4468: out<=1;
   4469: out<=0;
   4470: out<=0;
   4471: out<=1;
   4472: out<=0;
   4473: out<=1;
   4474: out<=0;
   4475: out<=1;
   4476: out<=0;
   4477: out<=0;
   4478: out<=1;
   4479: out<=1;
   4480: out<=1;
   4481: out<=1;
   4482: out<=0;
   4483: out<=0;
   4484: out<=1;
   4485: out<=0;
   4486: out<=1;
   4487: out<=0;
   4488: out<=1;
   4489: out<=0;
   4490: out<=0;
   4491: out<=1;
   4492: out<=1;
   4493: out<=1;
   4494: out<=1;
   4495: out<=1;
   4496: out<=0;
   4497: out<=1;
   4498: out<=0;
   4499: out<=1;
   4500: out<=1;
   4501: out<=1;
   4502: out<=0;
   4503: out<=0;
   4504: out<=1;
   4505: out<=1;
   4506: out<=1;
   4507: out<=1;
   4508: out<=0;
   4509: out<=1;
   4510: out<=1;
   4511: out<=0;
   4512: out<=0;
   4513: out<=1;
   4514: out<=1;
   4515: out<=0;
   4516: out<=1;
   4517: out<=1;
   4518: out<=1;
   4519: out<=1;
   4520: out<=0;
   4521: out<=0;
   4522: out<=1;
   4523: out<=1;
   4524: out<=1;
   4525: out<=0;
   4526: out<=1;
   4527: out<=0;
   4528: out<=1;
   4529: out<=1;
   4530: out<=1;
   4531: out<=1;
   4532: out<=1;
   4533: out<=0;
   4534: out<=0;
   4535: out<=1;
   4536: out<=0;
   4537: out<=1;
   4538: out<=0;
   4539: out<=1;
   4540: out<=0;
   4541: out<=0;
   4542: out<=1;
   4543: out<=1;
   4544: out<=1;
   4545: out<=1;
   4546: out<=0;
   4547: out<=0;
   4548: out<=1;
   4549: out<=0;
   4550: out<=1;
   4551: out<=0;
   4552: out<=1;
   4553: out<=0;
   4554: out<=0;
   4555: out<=1;
   4556: out<=1;
   4557: out<=1;
   4558: out<=1;
   4559: out<=1;
   4560: out<=1;
   4561: out<=0;
   4562: out<=1;
   4563: out<=0;
   4564: out<=0;
   4565: out<=0;
   4566: out<=1;
   4567: out<=1;
   4568: out<=0;
   4569: out<=0;
   4570: out<=0;
   4571: out<=0;
   4572: out<=1;
   4573: out<=0;
   4574: out<=0;
   4575: out<=1;
   4576: out<=1;
   4577: out<=0;
   4578: out<=0;
   4579: out<=1;
   4580: out<=0;
   4581: out<=0;
   4582: out<=0;
   4583: out<=0;
   4584: out<=1;
   4585: out<=1;
   4586: out<=0;
   4587: out<=0;
   4588: out<=0;
   4589: out<=1;
   4590: out<=0;
   4591: out<=1;
   4592: out<=1;
   4593: out<=1;
   4594: out<=1;
   4595: out<=1;
   4596: out<=1;
   4597: out<=0;
   4598: out<=0;
   4599: out<=1;
   4600: out<=0;
   4601: out<=1;
   4602: out<=0;
   4603: out<=1;
   4604: out<=0;
   4605: out<=0;
   4606: out<=1;
   4607: out<=1;
   4608: out<=1;
   4609: out<=1;
   4610: out<=1;
   4611: out<=1;
   4612: out<=1;
   4613: out<=0;
   4614: out<=0;
   4615: out<=1;
   4616: out<=0;
   4617: out<=1;
   4618: out<=0;
   4619: out<=1;
   4620: out<=0;
   4621: out<=0;
   4622: out<=1;
   4623: out<=1;
   4624: out<=1;
   4625: out<=0;
   4626: out<=0;
   4627: out<=1;
   4628: out<=0;
   4629: out<=0;
   4630: out<=0;
   4631: out<=0;
   4632: out<=1;
   4633: out<=1;
   4634: out<=0;
   4635: out<=0;
   4636: out<=0;
   4637: out<=1;
   4638: out<=0;
   4639: out<=1;
   4640: out<=1;
   4641: out<=0;
   4642: out<=1;
   4643: out<=0;
   4644: out<=0;
   4645: out<=0;
   4646: out<=1;
   4647: out<=1;
   4648: out<=0;
   4649: out<=0;
   4650: out<=0;
   4651: out<=0;
   4652: out<=1;
   4653: out<=0;
   4654: out<=0;
   4655: out<=1;
   4656: out<=1;
   4657: out<=1;
   4658: out<=0;
   4659: out<=0;
   4660: out<=1;
   4661: out<=0;
   4662: out<=1;
   4663: out<=0;
   4664: out<=1;
   4665: out<=0;
   4666: out<=0;
   4667: out<=1;
   4668: out<=1;
   4669: out<=1;
   4670: out<=1;
   4671: out<=1;
   4672: out<=1;
   4673: out<=1;
   4674: out<=1;
   4675: out<=1;
   4676: out<=1;
   4677: out<=0;
   4678: out<=0;
   4679: out<=1;
   4680: out<=0;
   4681: out<=1;
   4682: out<=0;
   4683: out<=1;
   4684: out<=0;
   4685: out<=0;
   4686: out<=1;
   4687: out<=1;
   4688: out<=0;
   4689: out<=1;
   4690: out<=1;
   4691: out<=0;
   4692: out<=1;
   4693: out<=1;
   4694: out<=1;
   4695: out<=1;
   4696: out<=0;
   4697: out<=0;
   4698: out<=1;
   4699: out<=1;
   4700: out<=1;
   4701: out<=0;
   4702: out<=1;
   4703: out<=0;
   4704: out<=0;
   4705: out<=1;
   4706: out<=0;
   4707: out<=1;
   4708: out<=1;
   4709: out<=1;
   4710: out<=0;
   4711: out<=0;
   4712: out<=1;
   4713: out<=1;
   4714: out<=1;
   4715: out<=1;
   4716: out<=0;
   4717: out<=1;
   4718: out<=1;
   4719: out<=0;
   4720: out<=1;
   4721: out<=1;
   4722: out<=0;
   4723: out<=0;
   4724: out<=1;
   4725: out<=0;
   4726: out<=1;
   4727: out<=0;
   4728: out<=1;
   4729: out<=0;
   4730: out<=0;
   4731: out<=1;
   4732: out<=1;
   4733: out<=1;
   4734: out<=1;
   4735: out<=1;
   4736: out<=1;
   4737: out<=1;
   4738: out<=1;
   4739: out<=1;
   4740: out<=1;
   4741: out<=0;
   4742: out<=0;
   4743: out<=1;
   4744: out<=0;
   4745: out<=1;
   4746: out<=0;
   4747: out<=1;
   4748: out<=0;
   4749: out<=0;
   4750: out<=1;
   4751: out<=1;
   4752: out<=0;
   4753: out<=1;
   4754: out<=1;
   4755: out<=0;
   4756: out<=1;
   4757: out<=1;
   4758: out<=1;
   4759: out<=1;
   4760: out<=0;
   4761: out<=0;
   4762: out<=1;
   4763: out<=1;
   4764: out<=1;
   4765: out<=0;
   4766: out<=1;
   4767: out<=0;
   4768: out<=1;
   4769: out<=0;
   4770: out<=1;
   4771: out<=0;
   4772: out<=0;
   4773: out<=0;
   4774: out<=1;
   4775: out<=1;
   4776: out<=0;
   4777: out<=0;
   4778: out<=0;
   4779: out<=0;
   4780: out<=1;
   4781: out<=0;
   4782: out<=0;
   4783: out<=1;
   4784: out<=0;
   4785: out<=0;
   4786: out<=1;
   4787: out<=1;
   4788: out<=0;
   4789: out<=1;
   4790: out<=0;
   4791: out<=1;
   4792: out<=0;
   4793: out<=1;
   4794: out<=1;
   4795: out<=0;
   4796: out<=0;
   4797: out<=0;
   4798: out<=0;
   4799: out<=0;
   4800: out<=1;
   4801: out<=1;
   4802: out<=1;
   4803: out<=1;
   4804: out<=1;
   4805: out<=0;
   4806: out<=0;
   4807: out<=1;
   4808: out<=0;
   4809: out<=1;
   4810: out<=0;
   4811: out<=1;
   4812: out<=0;
   4813: out<=0;
   4814: out<=1;
   4815: out<=1;
   4816: out<=1;
   4817: out<=0;
   4818: out<=0;
   4819: out<=1;
   4820: out<=0;
   4821: out<=0;
   4822: out<=0;
   4823: out<=0;
   4824: out<=1;
   4825: out<=1;
   4826: out<=0;
   4827: out<=0;
   4828: out<=0;
   4829: out<=1;
   4830: out<=0;
   4831: out<=1;
   4832: out<=0;
   4833: out<=1;
   4834: out<=0;
   4835: out<=1;
   4836: out<=1;
   4837: out<=1;
   4838: out<=0;
   4839: out<=0;
   4840: out<=1;
   4841: out<=1;
   4842: out<=1;
   4843: out<=1;
   4844: out<=0;
   4845: out<=1;
   4846: out<=1;
   4847: out<=0;
   4848: out<=0;
   4849: out<=0;
   4850: out<=1;
   4851: out<=1;
   4852: out<=0;
   4853: out<=1;
   4854: out<=0;
   4855: out<=1;
   4856: out<=0;
   4857: out<=1;
   4858: out<=1;
   4859: out<=0;
   4860: out<=0;
   4861: out<=0;
   4862: out<=0;
   4863: out<=0;
   4864: out<=0;
   4865: out<=1;
   4866: out<=1;
   4867: out<=0;
   4868: out<=1;
   4869: out<=1;
   4870: out<=1;
   4871: out<=1;
   4872: out<=0;
   4873: out<=0;
   4874: out<=1;
   4875: out<=1;
   4876: out<=1;
   4877: out<=0;
   4878: out<=1;
   4879: out<=0;
   4880: out<=1;
   4881: out<=1;
   4882: out<=1;
   4883: out<=1;
   4884: out<=1;
   4885: out<=0;
   4886: out<=0;
   4887: out<=1;
   4888: out<=0;
   4889: out<=1;
   4890: out<=0;
   4891: out<=1;
   4892: out<=0;
   4893: out<=0;
   4894: out<=1;
   4895: out<=1;
   4896: out<=1;
   4897: out<=1;
   4898: out<=0;
   4899: out<=0;
   4900: out<=1;
   4901: out<=0;
   4902: out<=1;
   4903: out<=0;
   4904: out<=1;
   4905: out<=0;
   4906: out<=0;
   4907: out<=1;
   4908: out<=1;
   4909: out<=1;
   4910: out<=1;
   4911: out<=1;
   4912: out<=0;
   4913: out<=1;
   4914: out<=0;
   4915: out<=1;
   4916: out<=1;
   4917: out<=1;
   4918: out<=0;
   4919: out<=0;
   4920: out<=1;
   4921: out<=1;
   4922: out<=1;
   4923: out<=1;
   4924: out<=0;
   4925: out<=1;
   4926: out<=1;
   4927: out<=0;
   4928: out<=1;
   4929: out<=0;
   4930: out<=0;
   4931: out<=1;
   4932: out<=0;
   4933: out<=0;
   4934: out<=0;
   4935: out<=0;
   4936: out<=1;
   4937: out<=1;
   4938: out<=0;
   4939: out<=0;
   4940: out<=0;
   4941: out<=1;
   4942: out<=0;
   4943: out<=1;
   4944: out<=1;
   4945: out<=1;
   4946: out<=1;
   4947: out<=1;
   4948: out<=1;
   4949: out<=0;
   4950: out<=0;
   4951: out<=1;
   4952: out<=0;
   4953: out<=1;
   4954: out<=0;
   4955: out<=1;
   4956: out<=0;
   4957: out<=0;
   4958: out<=1;
   4959: out<=1;
   4960: out<=1;
   4961: out<=1;
   4962: out<=0;
   4963: out<=0;
   4964: out<=1;
   4965: out<=0;
   4966: out<=1;
   4967: out<=0;
   4968: out<=1;
   4969: out<=0;
   4970: out<=0;
   4971: out<=1;
   4972: out<=1;
   4973: out<=1;
   4974: out<=1;
   4975: out<=1;
   4976: out<=1;
   4977: out<=0;
   4978: out<=1;
   4979: out<=0;
   4980: out<=0;
   4981: out<=0;
   4982: out<=1;
   4983: out<=1;
   4984: out<=0;
   4985: out<=0;
   4986: out<=0;
   4987: out<=0;
   4988: out<=1;
   4989: out<=0;
   4990: out<=0;
   4991: out<=1;
   4992: out<=1;
   4993: out<=0;
   4994: out<=0;
   4995: out<=1;
   4996: out<=0;
   4997: out<=0;
   4998: out<=0;
   4999: out<=0;
   5000: out<=1;
   5001: out<=1;
   5002: out<=0;
   5003: out<=0;
   5004: out<=0;
   5005: out<=1;
   5006: out<=0;
   5007: out<=1;
   5008: out<=1;
   5009: out<=1;
   5010: out<=1;
   5011: out<=1;
   5012: out<=1;
   5013: out<=0;
   5014: out<=0;
   5015: out<=1;
   5016: out<=0;
   5017: out<=1;
   5018: out<=0;
   5019: out<=1;
   5020: out<=0;
   5021: out<=0;
   5022: out<=1;
   5023: out<=1;
   5024: out<=0;
   5025: out<=0;
   5026: out<=1;
   5027: out<=1;
   5028: out<=0;
   5029: out<=1;
   5030: out<=0;
   5031: out<=1;
   5032: out<=0;
   5033: out<=1;
   5034: out<=1;
   5035: out<=0;
   5036: out<=0;
   5037: out<=0;
   5038: out<=0;
   5039: out<=0;
   5040: out<=0;
   5041: out<=1;
   5042: out<=0;
   5043: out<=1;
   5044: out<=1;
   5045: out<=1;
   5046: out<=0;
   5047: out<=0;
   5048: out<=1;
   5049: out<=1;
   5050: out<=1;
   5051: out<=1;
   5052: out<=0;
   5053: out<=1;
   5054: out<=1;
   5055: out<=0;
   5056: out<=0;
   5057: out<=1;
   5058: out<=1;
   5059: out<=0;
   5060: out<=1;
   5061: out<=1;
   5062: out<=1;
   5063: out<=1;
   5064: out<=0;
   5065: out<=0;
   5066: out<=1;
   5067: out<=1;
   5068: out<=1;
   5069: out<=0;
   5070: out<=1;
   5071: out<=0;
   5072: out<=1;
   5073: out<=1;
   5074: out<=1;
   5075: out<=1;
   5076: out<=1;
   5077: out<=0;
   5078: out<=0;
   5079: out<=1;
   5080: out<=0;
   5081: out<=1;
   5082: out<=0;
   5083: out<=1;
   5084: out<=0;
   5085: out<=0;
   5086: out<=1;
   5087: out<=1;
   5088: out<=0;
   5089: out<=0;
   5090: out<=1;
   5091: out<=1;
   5092: out<=0;
   5093: out<=1;
   5094: out<=0;
   5095: out<=1;
   5096: out<=0;
   5097: out<=1;
   5098: out<=1;
   5099: out<=0;
   5100: out<=0;
   5101: out<=0;
   5102: out<=0;
   5103: out<=0;
   5104: out<=1;
   5105: out<=0;
   5106: out<=1;
   5107: out<=0;
   5108: out<=0;
   5109: out<=0;
   5110: out<=1;
   5111: out<=1;
   5112: out<=0;
   5113: out<=0;
   5114: out<=0;
   5115: out<=0;
   5116: out<=1;
   5117: out<=0;
   5118: out<=0;
   5119: out<=1;
   5120: out<=0;
   5121: out<=0;
   5122: out<=1;
   5123: out<=1;
   5124: out<=1;
   5125: out<=0;
   5126: out<=1;
   5127: out<=0;
   5128: out<=1;
   5129: out<=0;
   5130: out<=0;
   5131: out<=1;
   5132: out<=0;
   5133: out<=0;
   5134: out<=0;
   5135: out<=0;
   5136: out<=1;
   5137: out<=0;
   5138: out<=1;
   5139: out<=0;
   5140: out<=1;
   5141: out<=1;
   5142: out<=0;
   5143: out<=0;
   5144: out<=1;
   5145: out<=1;
   5146: out<=1;
   5147: out<=1;
   5148: out<=1;
   5149: out<=0;
   5150: out<=0;
   5151: out<=1;
   5152: out<=0;
   5153: out<=1;
   5154: out<=1;
   5155: out<=0;
   5156: out<=0;
   5157: out<=0;
   5158: out<=0;
   5159: out<=0;
   5160: out<=1;
   5161: out<=1;
   5162: out<=0;
   5163: out<=0;
   5164: out<=1;
   5165: out<=0;
   5166: out<=1;
   5167: out<=0;
   5168: out<=1;
   5169: out<=1;
   5170: out<=1;
   5171: out<=1;
   5172: out<=0;
   5173: out<=1;
   5174: out<=1;
   5175: out<=0;
   5176: out<=1;
   5177: out<=0;
   5178: out<=1;
   5179: out<=0;
   5180: out<=0;
   5181: out<=0;
   5182: out<=1;
   5183: out<=1;
   5184: out<=0;
   5185: out<=0;
   5186: out<=1;
   5187: out<=1;
   5188: out<=1;
   5189: out<=0;
   5190: out<=1;
   5191: out<=0;
   5192: out<=1;
   5193: out<=0;
   5194: out<=0;
   5195: out<=1;
   5196: out<=0;
   5197: out<=0;
   5198: out<=0;
   5199: out<=0;
   5200: out<=0;
   5201: out<=1;
   5202: out<=0;
   5203: out<=1;
   5204: out<=0;
   5205: out<=0;
   5206: out<=1;
   5207: out<=1;
   5208: out<=0;
   5209: out<=0;
   5210: out<=0;
   5211: out<=0;
   5212: out<=0;
   5213: out<=1;
   5214: out<=1;
   5215: out<=0;
   5216: out<=1;
   5217: out<=0;
   5218: out<=0;
   5219: out<=1;
   5220: out<=1;
   5221: out<=1;
   5222: out<=1;
   5223: out<=1;
   5224: out<=0;
   5225: out<=0;
   5226: out<=1;
   5227: out<=1;
   5228: out<=0;
   5229: out<=1;
   5230: out<=0;
   5231: out<=1;
   5232: out<=1;
   5233: out<=1;
   5234: out<=1;
   5235: out<=1;
   5236: out<=0;
   5237: out<=1;
   5238: out<=1;
   5239: out<=0;
   5240: out<=1;
   5241: out<=0;
   5242: out<=1;
   5243: out<=0;
   5244: out<=0;
   5245: out<=0;
   5246: out<=1;
   5247: out<=1;
   5248: out<=1;
   5249: out<=1;
   5250: out<=0;
   5251: out<=0;
   5252: out<=0;
   5253: out<=1;
   5254: out<=0;
   5255: out<=1;
   5256: out<=0;
   5257: out<=1;
   5258: out<=1;
   5259: out<=0;
   5260: out<=1;
   5261: out<=1;
   5262: out<=1;
   5263: out<=1;
   5264: out<=1;
   5265: out<=0;
   5266: out<=1;
   5267: out<=0;
   5268: out<=1;
   5269: out<=1;
   5270: out<=0;
   5271: out<=0;
   5272: out<=1;
   5273: out<=1;
   5274: out<=1;
   5275: out<=1;
   5276: out<=1;
   5277: out<=0;
   5278: out<=0;
   5279: out<=1;
   5280: out<=1;
   5281: out<=0;
   5282: out<=0;
   5283: out<=1;
   5284: out<=1;
   5285: out<=1;
   5286: out<=1;
   5287: out<=1;
   5288: out<=0;
   5289: out<=0;
   5290: out<=1;
   5291: out<=1;
   5292: out<=0;
   5293: out<=1;
   5294: out<=0;
   5295: out<=1;
   5296: out<=1;
   5297: out<=1;
   5298: out<=1;
   5299: out<=1;
   5300: out<=0;
   5301: out<=1;
   5302: out<=1;
   5303: out<=0;
   5304: out<=1;
   5305: out<=0;
   5306: out<=1;
   5307: out<=0;
   5308: out<=0;
   5309: out<=0;
   5310: out<=1;
   5311: out<=1;
   5312: out<=1;
   5313: out<=1;
   5314: out<=0;
   5315: out<=0;
   5316: out<=0;
   5317: out<=1;
   5318: out<=0;
   5319: out<=1;
   5320: out<=0;
   5321: out<=1;
   5322: out<=1;
   5323: out<=0;
   5324: out<=1;
   5325: out<=1;
   5326: out<=1;
   5327: out<=1;
   5328: out<=0;
   5329: out<=1;
   5330: out<=0;
   5331: out<=1;
   5332: out<=0;
   5333: out<=0;
   5334: out<=1;
   5335: out<=1;
   5336: out<=0;
   5337: out<=0;
   5338: out<=0;
   5339: out<=0;
   5340: out<=0;
   5341: out<=1;
   5342: out<=1;
   5343: out<=0;
   5344: out<=0;
   5345: out<=1;
   5346: out<=1;
   5347: out<=0;
   5348: out<=0;
   5349: out<=0;
   5350: out<=0;
   5351: out<=0;
   5352: out<=1;
   5353: out<=1;
   5354: out<=0;
   5355: out<=0;
   5356: out<=1;
   5357: out<=0;
   5358: out<=1;
   5359: out<=0;
   5360: out<=1;
   5361: out<=1;
   5362: out<=1;
   5363: out<=1;
   5364: out<=0;
   5365: out<=1;
   5366: out<=1;
   5367: out<=0;
   5368: out<=1;
   5369: out<=0;
   5370: out<=1;
   5371: out<=0;
   5372: out<=0;
   5373: out<=0;
   5374: out<=1;
   5375: out<=1;
   5376: out<=0;
   5377: out<=1;
   5378: out<=0;
   5379: out<=1;
   5380: out<=0;
   5381: out<=0;
   5382: out<=1;
   5383: out<=1;
   5384: out<=0;
   5385: out<=0;
   5386: out<=0;
   5387: out<=0;
   5388: out<=0;
   5389: out<=1;
   5390: out<=1;
   5391: out<=0;
   5392: out<=0;
   5393: out<=0;
   5394: out<=1;
   5395: out<=1;
   5396: out<=1;
   5397: out<=0;
   5398: out<=1;
   5399: out<=0;
   5400: out<=1;
   5401: out<=0;
   5402: out<=0;
   5403: out<=1;
   5404: out<=0;
   5405: out<=0;
   5406: out<=0;
   5407: out<=0;
   5408: out<=1;
   5409: out<=1;
   5410: out<=1;
   5411: out<=1;
   5412: out<=0;
   5413: out<=1;
   5414: out<=1;
   5415: out<=0;
   5416: out<=1;
   5417: out<=0;
   5418: out<=1;
   5419: out<=0;
   5420: out<=0;
   5421: out<=0;
   5422: out<=1;
   5423: out<=1;
   5424: out<=1;
   5425: out<=0;
   5426: out<=0;
   5427: out<=1;
   5428: out<=1;
   5429: out<=1;
   5430: out<=1;
   5431: out<=1;
   5432: out<=0;
   5433: out<=0;
   5434: out<=1;
   5435: out<=1;
   5436: out<=0;
   5437: out<=1;
   5438: out<=0;
   5439: out<=1;
   5440: out<=1;
   5441: out<=0;
   5442: out<=1;
   5443: out<=0;
   5444: out<=1;
   5445: out<=1;
   5446: out<=0;
   5447: out<=0;
   5448: out<=1;
   5449: out<=1;
   5450: out<=1;
   5451: out<=1;
   5452: out<=1;
   5453: out<=0;
   5454: out<=0;
   5455: out<=1;
   5456: out<=0;
   5457: out<=0;
   5458: out<=1;
   5459: out<=1;
   5460: out<=1;
   5461: out<=0;
   5462: out<=1;
   5463: out<=0;
   5464: out<=1;
   5465: out<=0;
   5466: out<=0;
   5467: out<=1;
   5468: out<=0;
   5469: out<=0;
   5470: out<=0;
   5471: out<=0;
   5472: out<=1;
   5473: out<=1;
   5474: out<=1;
   5475: out<=1;
   5476: out<=0;
   5477: out<=1;
   5478: out<=1;
   5479: out<=0;
   5480: out<=1;
   5481: out<=0;
   5482: out<=1;
   5483: out<=0;
   5484: out<=0;
   5485: out<=0;
   5486: out<=1;
   5487: out<=1;
   5488: out<=0;
   5489: out<=1;
   5490: out<=1;
   5491: out<=0;
   5492: out<=0;
   5493: out<=0;
   5494: out<=0;
   5495: out<=0;
   5496: out<=1;
   5497: out<=1;
   5498: out<=0;
   5499: out<=0;
   5500: out<=1;
   5501: out<=0;
   5502: out<=1;
   5503: out<=0;
   5504: out<=0;
   5505: out<=1;
   5506: out<=0;
   5507: out<=1;
   5508: out<=0;
   5509: out<=0;
   5510: out<=1;
   5511: out<=1;
   5512: out<=0;
   5513: out<=0;
   5514: out<=0;
   5515: out<=0;
   5516: out<=0;
   5517: out<=1;
   5518: out<=1;
   5519: out<=0;
   5520: out<=1;
   5521: out<=1;
   5522: out<=0;
   5523: out<=0;
   5524: out<=0;
   5525: out<=1;
   5526: out<=0;
   5527: out<=1;
   5528: out<=0;
   5529: out<=1;
   5530: out<=1;
   5531: out<=0;
   5532: out<=1;
   5533: out<=1;
   5534: out<=1;
   5535: out<=1;
   5536: out<=1;
   5537: out<=1;
   5538: out<=1;
   5539: out<=1;
   5540: out<=0;
   5541: out<=1;
   5542: out<=1;
   5543: out<=0;
   5544: out<=1;
   5545: out<=0;
   5546: out<=1;
   5547: out<=0;
   5548: out<=0;
   5549: out<=0;
   5550: out<=1;
   5551: out<=1;
   5552: out<=0;
   5553: out<=1;
   5554: out<=1;
   5555: out<=0;
   5556: out<=0;
   5557: out<=0;
   5558: out<=0;
   5559: out<=0;
   5560: out<=1;
   5561: out<=1;
   5562: out<=0;
   5563: out<=0;
   5564: out<=1;
   5565: out<=0;
   5566: out<=1;
   5567: out<=0;
   5568: out<=1;
   5569: out<=0;
   5570: out<=1;
   5571: out<=0;
   5572: out<=1;
   5573: out<=1;
   5574: out<=0;
   5575: out<=0;
   5576: out<=1;
   5577: out<=1;
   5578: out<=1;
   5579: out<=1;
   5580: out<=1;
   5581: out<=0;
   5582: out<=0;
   5583: out<=1;
   5584: out<=1;
   5585: out<=1;
   5586: out<=0;
   5587: out<=0;
   5588: out<=0;
   5589: out<=1;
   5590: out<=0;
   5591: out<=1;
   5592: out<=0;
   5593: out<=1;
   5594: out<=1;
   5595: out<=0;
   5596: out<=1;
   5597: out<=1;
   5598: out<=1;
   5599: out<=1;
   5600: out<=1;
   5601: out<=1;
   5602: out<=1;
   5603: out<=1;
   5604: out<=0;
   5605: out<=1;
   5606: out<=1;
   5607: out<=0;
   5608: out<=1;
   5609: out<=0;
   5610: out<=1;
   5611: out<=0;
   5612: out<=0;
   5613: out<=0;
   5614: out<=1;
   5615: out<=1;
   5616: out<=1;
   5617: out<=0;
   5618: out<=0;
   5619: out<=1;
   5620: out<=1;
   5621: out<=1;
   5622: out<=1;
   5623: out<=1;
   5624: out<=0;
   5625: out<=0;
   5626: out<=1;
   5627: out<=1;
   5628: out<=0;
   5629: out<=1;
   5630: out<=0;
   5631: out<=1;
   5632: out<=1;
   5633: out<=0;
   5634: out<=0;
   5635: out<=1;
   5636: out<=1;
   5637: out<=1;
   5638: out<=1;
   5639: out<=1;
   5640: out<=0;
   5641: out<=0;
   5642: out<=1;
   5643: out<=1;
   5644: out<=0;
   5645: out<=1;
   5646: out<=0;
   5647: out<=1;
   5648: out<=1;
   5649: out<=1;
   5650: out<=1;
   5651: out<=1;
   5652: out<=0;
   5653: out<=1;
   5654: out<=1;
   5655: out<=0;
   5656: out<=1;
   5657: out<=0;
   5658: out<=1;
   5659: out<=0;
   5660: out<=0;
   5661: out<=0;
   5662: out<=1;
   5663: out<=1;
   5664: out<=1;
   5665: out<=1;
   5666: out<=0;
   5667: out<=0;
   5668: out<=0;
   5669: out<=1;
   5670: out<=0;
   5671: out<=1;
   5672: out<=0;
   5673: out<=1;
   5674: out<=1;
   5675: out<=0;
   5676: out<=1;
   5677: out<=1;
   5678: out<=1;
   5679: out<=1;
   5680: out<=1;
   5681: out<=0;
   5682: out<=1;
   5683: out<=0;
   5684: out<=1;
   5685: out<=1;
   5686: out<=0;
   5687: out<=0;
   5688: out<=1;
   5689: out<=1;
   5690: out<=1;
   5691: out<=1;
   5692: out<=1;
   5693: out<=0;
   5694: out<=0;
   5695: out<=1;
   5696: out<=0;
   5697: out<=1;
   5698: out<=1;
   5699: out<=0;
   5700: out<=0;
   5701: out<=0;
   5702: out<=0;
   5703: out<=0;
   5704: out<=1;
   5705: out<=1;
   5706: out<=0;
   5707: out<=0;
   5708: out<=1;
   5709: out<=0;
   5710: out<=1;
   5711: out<=0;
   5712: out<=1;
   5713: out<=1;
   5714: out<=1;
   5715: out<=1;
   5716: out<=0;
   5717: out<=1;
   5718: out<=1;
   5719: out<=0;
   5720: out<=1;
   5721: out<=0;
   5722: out<=1;
   5723: out<=0;
   5724: out<=0;
   5725: out<=0;
   5726: out<=1;
   5727: out<=1;
   5728: out<=1;
   5729: out<=1;
   5730: out<=0;
   5731: out<=0;
   5732: out<=0;
   5733: out<=1;
   5734: out<=0;
   5735: out<=1;
   5736: out<=0;
   5737: out<=1;
   5738: out<=1;
   5739: out<=0;
   5740: out<=1;
   5741: out<=1;
   5742: out<=1;
   5743: out<=1;
   5744: out<=0;
   5745: out<=1;
   5746: out<=0;
   5747: out<=1;
   5748: out<=0;
   5749: out<=0;
   5750: out<=1;
   5751: out<=1;
   5752: out<=0;
   5753: out<=0;
   5754: out<=0;
   5755: out<=0;
   5756: out<=0;
   5757: out<=1;
   5758: out<=1;
   5759: out<=0;
   5760: out<=0;
   5761: out<=1;
   5762: out<=1;
   5763: out<=0;
   5764: out<=0;
   5765: out<=0;
   5766: out<=0;
   5767: out<=0;
   5768: out<=1;
   5769: out<=1;
   5770: out<=0;
   5771: out<=0;
   5772: out<=1;
   5773: out<=0;
   5774: out<=1;
   5775: out<=0;
   5776: out<=1;
   5777: out<=1;
   5778: out<=1;
   5779: out<=1;
   5780: out<=0;
   5781: out<=1;
   5782: out<=1;
   5783: out<=0;
   5784: out<=1;
   5785: out<=0;
   5786: out<=1;
   5787: out<=0;
   5788: out<=0;
   5789: out<=0;
   5790: out<=1;
   5791: out<=1;
   5792: out<=0;
   5793: out<=0;
   5794: out<=1;
   5795: out<=1;
   5796: out<=1;
   5797: out<=0;
   5798: out<=1;
   5799: out<=0;
   5800: out<=1;
   5801: out<=0;
   5802: out<=0;
   5803: out<=1;
   5804: out<=0;
   5805: out<=0;
   5806: out<=0;
   5807: out<=0;
   5808: out<=1;
   5809: out<=0;
   5810: out<=1;
   5811: out<=0;
   5812: out<=1;
   5813: out<=1;
   5814: out<=0;
   5815: out<=0;
   5816: out<=1;
   5817: out<=1;
   5818: out<=1;
   5819: out<=1;
   5820: out<=1;
   5821: out<=0;
   5822: out<=0;
   5823: out<=1;
   5824: out<=1;
   5825: out<=0;
   5826: out<=0;
   5827: out<=1;
   5828: out<=1;
   5829: out<=1;
   5830: out<=1;
   5831: out<=1;
   5832: out<=0;
   5833: out<=0;
   5834: out<=1;
   5835: out<=1;
   5836: out<=0;
   5837: out<=1;
   5838: out<=0;
   5839: out<=1;
   5840: out<=1;
   5841: out<=1;
   5842: out<=1;
   5843: out<=1;
   5844: out<=0;
   5845: out<=1;
   5846: out<=1;
   5847: out<=0;
   5848: out<=1;
   5849: out<=0;
   5850: out<=1;
   5851: out<=0;
   5852: out<=0;
   5853: out<=0;
   5854: out<=1;
   5855: out<=1;
   5856: out<=0;
   5857: out<=0;
   5858: out<=1;
   5859: out<=1;
   5860: out<=1;
   5861: out<=0;
   5862: out<=1;
   5863: out<=0;
   5864: out<=1;
   5865: out<=0;
   5866: out<=0;
   5867: out<=1;
   5868: out<=0;
   5869: out<=0;
   5870: out<=0;
   5871: out<=0;
   5872: out<=0;
   5873: out<=1;
   5874: out<=0;
   5875: out<=1;
   5876: out<=0;
   5877: out<=0;
   5878: out<=1;
   5879: out<=1;
   5880: out<=0;
   5881: out<=0;
   5882: out<=0;
   5883: out<=0;
   5884: out<=0;
   5885: out<=1;
   5886: out<=1;
   5887: out<=0;
   5888: out<=1;
   5889: out<=1;
   5890: out<=1;
   5891: out<=1;
   5892: out<=0;
   5893: out<=1;
   5894: out<=1;
   5895: out<=0;
   5896: out<=1;
   5897: out<=0;
   5898: out<=1;
   5899: out<=0;
   5900: out<=0;
   5901: out<=0;
   5902: out<=1;
   5903: out<=1;
   5904: out<=0;
   5905: out<=1;
   5906: out<=1;
   5907: out<=0;
   5908: out<=0;
   5909: out<=0;
   5910: out<=0;
   5911: out<=0;
   5912: out<=1;
   5913: out<=1;
   5914: out<=0;
   5915: out<=0;
   5916: out<=1;
   5917: out<=0;
   5918: out<=1;
   5919: out<=0;
   5920: out<=0;
   5921: out<=1;
   5922: out<=0;
   5923: out<=1;
   5924: out<=0;
   5925: out<=0;
   5926: out<=1;
   5927: out<=1;
   5928: out<=0;
   5929: out<=0;
   5930: out<=0;
   5931: out<=0;
   5932: out<=0;
   5933: out<=1;
   5934: out<=1;
   5935: out<=0;
   5936: out<=1;
   5937: out<=1;
   5938: out<=0;
   5939: out<=0;
   5940: out<=0;
   5941: out<=1;
   5942: out<=0;
   5943: out<=1;
   5944: out<=0;
   5945: out<=1;
   5946: out<=1;
   5947: out<=0;
   5948: out<=1;
   5949: out<=1;
   5950: out<=1;
   5951: out<=1;
   5952: out<=1;
   5953: out<=1;
   5954: out<=1;
   5955: out<=1;
   5956: out<=0;
   5957: out<=1;
   5958: out<=1;
   5959: out<=0;
   5960: out<=1;
   5961: out<=0;
   5962: out<=1;
   5963: out<=0;
   5964: out<=0;
   5965: out<=0;
   5966: out<=1;
   5967: out<=1;
   5968: out<=1;
   5969: out<=0;
   5970: out<=0;
   5971: out<=1;
   5972: out<=1;
   5973: out<=1;
   5974: out<=1;
   5975: out<=1;
   5976: out<=0;
   5977: out<=0;
   5978: out<=1;
   5979: out<=1;
   5980: out<=0;
   5981: out<=1;
   5982: out<=0;
   5983: out<=1;
   5984: out<=1;
   5985: out<=0;
   5986: out<=1;
   5987: out<=0;
   5988: out<=1;
   5989: out<=1;
   5990: out<=0;
   5991: out<=0;
   5992: out<=1;
   5993: out<=1;
   5994: out<=1;
   5995: out<=1;
   5996: out<=1;
   5997: out<=0;
   5998: out<=0;
   5999: out<=1;
   6000: out<=1;
   6001: out<=1;
   6002: out<=0;
   6003: out<=0;
   6004: out<=0;
   6005: out<=1;
   6006: out<=0;
   6007: out<=1;
   6008: out<=0;
   6009: out<=1;
   6010: out<=1;
   6011: out<=0;
   6012: out<=1;
   6013: out<=1;
   6014: out<=1;
   6015: out<=1;
   6016: out<=1;
   6017: out<=1;
   6018: out<=1;
   6019: out<=1;
   6020: out<=0;
   6021: out<=1;
   6022: out<=1;
   6023: out<=0;
   6024: out<=1;
   6025: out<=0;
   6026: out<=1;
   6027: out<=0;
   6028: out<=0;
   6029: out<=0;
   6030: out<=1;
   6031: out<=1;
   6032: out<=1;
   6033: out<=0;
   6034: out<=0;
   6035: out<=1;
   6036: out<=1;
   6037: out<=1;
   6038: out<=1;
   6039: out<=1;
   6040: out<=0;
   6041: out<=0;
   6042: out<=1;
   6043: out<=1;
   6044: out<=0;
   6045: out<=1;
   6046: out<=0;
   6047: out<=1;
   6048: out<=0;
   6049: out<=1;
   6050: out<=0;
   6051: out<=1;
   6052: out<=0;
   6053: out<=0;
   6054: out<=1;
   6055: out<=1;
   6056: out<=0;
   6057: out<=0;
   6058: out<=0;
   6059: out<=0;
   6060: out<=0;
   6061: out<=1;
   6062: out<=1;
   6063: out<=0;
   6064: out<=0;
   6065: out<=0;
   6066: out<=1;
   6067: out<=1;
   6068: out<=1;
   6069: out<=0;
   6070: out<=1;
   6071: out<=0;
   6072: out<=1;
   6073: out<=0;
   6074: out<=0;
   6075: out<=1;
   6076: out<=0;
   6077: out<=0;
   6078: out<=0;
   6079: out<=0;
   6080: out<=1;
   6081: out<=1;
   6082: out<=1;
   6083: out<=1;
   6084: out<=0;
   6085: out<=1;
   6086: out<=1;
   6087: out<=0;
   6088: out<=1;
   6089: out<=0;
   6090: out<=1;
   6091: out<=0;
   6092: out<=0;
   6093: out<=0;
   6094: out<=1;
   6095: out<=1;
   6096: out<=0;
   6097: out<=1;
   6098: out<=1;
   6099: out<=0;
   6100: out<=0;
   6101: out<=0;
   6102: out<=0;
   6103: out<=0;
   6104: out<=1;
   6105: out<=1;
   6106: out<=0;
   6107: out<=0;
   6108: out<=1;
   6109: out<=0;
   6110: out<=1;
   6111: out<=0;
   6112: out<=1;
   6113: out<=0;
   6114: out<=1;
   6115: out<=0;
   6116: out<=1;
   6117: out<=1;
   6118: out<=0;
   6119: out<=0;
   6120: out<=1;
   6121: out<=1;
   6122: out<=1;
   6123: out<=1;
   6124: out<=1;
   6125: out<=0;
   6126: out<=0;
   6127: out<=1;
   6128: out<=0;
   6129: out<=0;
   6130: out<=1;
   6131: out<=1;
   6132: out<=1;
   6133: out<=0;
   6134: out<=1;
   6135: out<=0;
   6136: out<=1;
   6137: out<=0;
   6138: out<=0;
   6139: out<=1;
   6140: out<=0;
   6141: out<=0;
   6142: out<=0;
   6143: out<=0;
   6144: out<=1;
   6145: out<=1;
   6146: out<=1;
   6147: out<=1;
   6148: out<=0;
   6149: out<=1;
   6150: out<=1;
   6151: out<=0;
   6152: out<=0;
   6153: out<=1;
   6154: out<=0;
   6155: out<=1;
   6156: out<=1;
   6157: out<=1;
   6158: out<=0;
   6159: out<=0;
   6160: out<=0;
   6161: out<=1;
   6162: out<=1;
   6163: out<=0;
   6164: out<=0;
   6165: out<=0;
   6166: out<=0;
   6167: out<=0;
   6168: out<=0;
   6169: out<=0;
   6170: out<=1;
   6171: out<=1;
   6172: out<=0;
   6173: out<=1;
   6174: out<=0;
   6175: out<=1;
   6176: out<=1;
   6177: out<=0;
   6178: out<=1;
   6179: out<=0;
   6180: out<=1;
   6181: out<=1;
   6182: out<=0;
   6183: out<=0;
   6184: out<=0;
   6185: out<=0;
   6186: out<=0;
   6187: out<=0;
   6188: out<=0;
   6189: out<=1;
   6190: out<=1;
   6191: out<=0;
   6192: out<=0;
   6193: out<=0;
   6194: out<=1;
   6195: out<=1;
   6196: out<=1;
   6197: out<=0;
   6198: out<=1;
   6199: out<=0;
   6200: out<=0;
   6201: out<=1;
   6202: out<=1;
   6203: out<=0;
   6204: out<=1;
   6205: out<=1;
   6206: out<=1;
   6207: out<=1;
   6208: out<=1;
   6209: out<=1;
   6210: out<=1;
   6211: out<=1;
   6212: out<=0;
   6213: out<=1;
   6214: out<=1;
   6215: out<=0;
   6216: out<=0;
   6217: out<=1;
   6218: out<=0;
   6219: out<=1;
   6220: out<=1;
   6221: out<=1;
   6222: out<=0;
   6223: out<=0;
   6224: out<=1;
   6225: out<=0;
   6226: out<=0;
   6227: out<=1;
   6228: out<=1;
   6229: out<=1;
   6230: out<=1;
   6231: out<=1;
   6232: out<=1;
   6233: out<=1;
   6234: out<=0;
   6235: out<=0;
   6236: out<=1;
   6237: out<=0;
   6238: out<=1;
   6239: out<=0;
   6240: out<=0;
   6241: out<=1;
   6242: out<=0;
   6243: out<=1;
   6244: out<=0;
   6245: out<=0;
   6246: out<=1;
   6247: out<=1;
   6248: out<=1;
   6249: out<=1;
   6250: out<=1;
   6251: out<=1;
   6252: out<=1;
   6253: out<=0;
   6254: out<=0;
   6255: out<=1;
   6256: out<=0;
   6257: out<=0;
   6258: out<=1;
   6259: out<=1;
   6260: out<=1;
   6261: out<=0;
   6262: out<=1;
   6263: out<=0;
   6264: out<=0;
   6265: out<=1;
   6266: out<=1;
   6267: out<=0;
   6268: out<=1;
   6269: out<=1;
   6270: out<=1;
   6271: out<=1;
   6272: out<=1;
   6273: out<=1;
   6274: out<=1;
   6275: out<=1;
   6276: out<=0;
   6277: out<=1;
   6278: out<=1;
   6279: out<=0;
   6280: out<=0;
   6281: out<=1;
   6282: out<=0;
   6283: out<=1;
   6284: out<=1;
   6285: out<=1;
   6286: out<=0;
   6287: out<=0;
   6288: out<=1;
   6289: out<=0;
   6290: out<=0;
   6291: out<=1;
   6292: out<=1;
   6293: out<=1;
   6294: out<=1;
   6295: out<=1;
   6296: out<=1;
   6297: out<=1;
   6298: out<=0;
   6299: out<=0;
   6300: out<=1;
   6301: out<=0;
   6302: out<=1;
   6303: out<=0;
   6304: out<=1;
   6305: out<=0;
   6306: out<=1;
   6307: out<=0;
   6308: out<=1;
   6309: out<=1;
   6310: out<=0;
   6311: out<=0;
   6312: out<=0;
   6313: out<=0;
   6314: out<=0;
   6315: out<=0;
   6316: out<=0;
   6317: out<=1;
   6318: out<=1;
   6319: out<=0;
   6320: out<=1;
   6321: out<=1;
   6322: out<=0;
   6323: out<=0;
   6324: out<=0;
   6325: out<=1;
   6326: out<=0;
   6327: out<=1;
   6328: out<=1;
   6329: out<=0;
   6330: out<=0;
   6331: out<=1;
   6332: out<=0;
   6333: out<=0;
   6334: out<=0;
   6335: out<=0;
   6336: out<=1;
   6337: out<=1;
   6338: out<=1;
   6339: out<=1;
   6340: out<=0;
   6341: out<=1;
   6342: out<=1;
   6343: out<=0;
   6344: out<=0;
   6345: out<=1;
   6346: out<=0;
   6347: out<=1;
   6348: out<=1;
   6349: out<=1;
   6350: out<=0;
   6351: out<=0;
   6352: out<=0;
   6353: out<=1;
   6354: out<=1;
   6355: out<=0;
   6356: out<=0;
   6357: out<=0;
   6358: out<=0;
   6359: out<=0;
   6360: out<=0;
   6361: out<=0;
   6362: out<=1;
   6363: out<=1;
   6364: out<=0;
   6365: out<=1;
   6366: out<=0;
   6367: out<=1;
   6368: out<=0;
   6369: out<=1;
   6370: out<=0;
   6371: out<=1;
   6372: out<=0;
   6373: out<=0;
   6374: out<=1;
   6375: out<=1;
   6376: out<=1;
   6377: out<=1;
   6378: out<=1;
   6379: out<=1;
   6380: out<=1;
   6381: out<=0;
   6382: out<=0;
   6383: out<=1;
   6384: out<=1;
   6385: out<=1;
   6386: out<=0;
   6387: out<=0;
   6388: out<=0;
   6389: out<=1;
   6390: out<=0;
   6391: out<=1;
   6392: out<=1;
   6393: out<=0;
   6394: out<=0;
   6395: out<=1;
   6396: out<=0;
   6397: out<=0;
   6398: out<=0;
   6399: out<=0;
   6400: out<=1;
   6401: out<=0;
   6402: out<=0;
   6403: out<=1;
   6404: out<=1;
   6405: out<=1;
   6406: out<=1;
   6407: out<=1;
   6408: out<=1;
   6409: out<=1;
   6410: out<=0;
   6411: out<=0;
   6412: out<=1;
   6413: out<=0;
   6414: out<=1;
   6415: out<=0;
   6416: out<=1;
   6417: out<=1;
   6418: out<=1;
   6419: out<=1;
   6420: out<=0;
   6421: out<=1;
   6422: out<=1;
   6423: out<=0;
   6424: out<=0;
   6425: out<=1;
   6426: out<=0;
   6427: out<=1;
   6428: out<=1;
   6429: out<=1;
   6430: out<=0;
   6431: out<=0;
   6432: out<=0;
   6433: out<=0;
   6434: out<=1;
   6435: out<=1;
   6436: out<=1;
   6437: out<=0;
   6438: out<=1;
   6439: out<=0;
   6440: out<=0;
   6441: out<=1;
   6442: out<=1;
   6443: out<=0;
   6444: out<=1;
   6445: out<=1;
   6446: out<=1;
   6447: out<=1;
   6448: out<=0;
   6449: out<=1;
   6450: out<=0;
   6451: out<=1;
   6452: out<=0;
   6453: out<=0;
   6454: out<=1;
   6455: out<=1;
   6456: out<=1;
   6457: out<=1;
   6458: out<=1;
   6459: out<=1;
   6460: out<=1;
   6461: out<=0;
   6462: out<=0;
   6463: out<=1;
   6464: out<=0;
   6465: out<=1;
   6466: out<=1;
   6467: out<=0;
   6468: out<=0;
   6469: out<=0;
   6470: out<=0;
   6471: out<=0;
   6472: out<=0;
   6473: out<=0;
   6474: out<=1;
   6475: out<=1;
   6476: out<=0;
   6477: out<=1;
   6478: out<=0;
   6479: out<=1;
   6480: out<=1;
   6481: out<=1;
   6482: out<=1;
   6483: out<=1;
   6484: out<=0;
   6485: out<=1;
   6486: out<=1;
   6487: out<=0;
   6488: out<=0;
   6489: out<=1;
   6490: out<=0;
   6491: out<=1;
   6492: out<=1;
   6493: out<=1;
   6494: out<=0;
   6495: out<=0;
   6496: out<=0;
   6497: out<=0;
   6498: out<=1;
   6499: out<=1;
   6500: out<=1;
   6501: out<=0;
   6502: out<=1;
   6503: out<=0;
   6504: out<=0;
   6505: out<=1;
   6506: out<=1;
   6507: out<=0;
   6508: out<=1;
   6509: out<=1;
   6510: out<=1;
   6511: out<=1;
   6512: out<=1;
   6513: out<=0;
   6514: out<=1;
   6515: out<=0;
   6516: out<=1;
   6517: out<=1;
   6518: out<=0;
   6519: out<=0;
   6520: out<=0;
   6521: out<=0;
   6522: out<=0;
   6523: out<=0;
   6524: out<=0;
   6525: out<=1;
   6526: out<=1;
   6527: out<=0;
   6528: out<=0;
   6529: out<=1;
   6530: out<=1;
   6531: out<=0;
   6532: out<=0;
   6533: out<=0;
   6534: out<=0;
   6535: out<=0;
   6536: out<=0;
   6537: out<=0;
   6538: out<=1;
   6539: out<=1;
   6540: out<=0;
   6541: out<=1;
   6542: out<=0;
   6543: out<=1;
   6544: out<=1;
   6545: out<=1;
   6546: out<=1;
   6547: out<=1;
   6548: out<=0;
   6549: out<=1;
   6550: out<=1;
   6551: out<=0;
   6552: out<=0;
   6553: out<=1;
   6554: out<=0;
   6555: out<=1;
   6556: out<=1;
   6557: out<=1;
   6558: out<=0;
   6559: out<=0;
   6560: out<=1;
   6561: out<=1;
   6562: out<=0;
   6563: out<=0;
   6564: out<=0;
   6565: out<=1;
   6566: out<=0;
   6567: out<=1;
   6568: out<=1;
   6569: out<=0;
   6570: out<=0;
   6571: out<=1;
   6572: out<=0;
   6573: out<=0;
   6574: out<=0;
   6575: out<=0;
   6576: out<=0;
   6577: out<=1;
   6578: out<=0;
   6579: out<=1;
   6580: out<=0;
   6581: out<=0;
   6582: out<=1;
   6583: out<=1;
   6584: out<=1;
   6585: out<=1;
   6586: out<=1;
   6587: out<=1;
   6588: out<=1;
   6589: out<=0;
   6590: out<=0;
   6591: out<=1;
   6592: out<=1;
   6593: out<=0;
   6594: out<=0;
   6595: out<=1;
   6596: out<=1;
   6597: out<=1;
   6598: out<=1;
   6599: out<=1;
   6600: out<=1;
   6601: out<=1;
   6602: out<=0;
   6603: out<=0;
   6604: out<=1;
   6605: out<=0;
   6606: out<=1;
   6607: out<=0;
   6608: out<=1;
   6609: out<=1;
   6610: out<=1;
   6611: out<=1;
   6612: out<=0;
   6613: out<=1;
   6614: out<=1;
   6615: out<=0;
   6616: out<=0;
   6617: out<=1;
   6618: out<=0;
   6619: out<=1;
   6620: out<=1;
   6621: out<=1;
   6622: out<=0;
   6623: out<=0;
   6624: out<=1;
   6625: out<=1;
   6626: out<=0;
   6627: out<=0;
   6628: out<=0;
   6629: out<=1;
   6630: out<=0;
   6631: out<=1;
   6632: out<=1;
   6633: out<=0;
   6634: out<=0;
   6635: out<=1;
   6636: out<=0;
   6637: out<=0;
   6638: out<=0;
   6639: out<=0;
   6640: out<=1;
   6641: out<=0;
   6642: out<=1;
   6643: out<=0;
   6644: out<=1;
   6645: out<=1;
   6646: out<=0;
   6647: out<=0;
   6648: out<=0;
   6649: out<=0;
   6650: out<=0;
   6651: out<=0;
   6652: out<=0;
   6653: out<=1;
   6654: out<=1;
   6655: out<=0;
   6656: out<=1;
   6657: out<=0;
   6658: out<=1;
   6659: out<=0;
   6660: out<=1;
   6661: out<=1;
   6662: out<=0;
   6663: out<=0;
   6664: out<=0;
   6665: out<=0;
   6666: out<=0;
   6667: out<=0;
   6668: out<=0;
   6669: out<=1;
   6670: out<=1;
   6671: out<=0;
   6672: out<=1;
   6673: out<=1;
   6674: out<=0;
   6675: out<=0;
   6676: out<=0;
   6677: out<=1;
   6678: out<=0;
   6679: out<=1;
   6680: out<=1;
   6681: out<=0;
   6682: out<=0;
   6683: out<=1;
   6684: out<=0;
   6685: out<=0;
   6686: out<=0;
   6687: out<=0;
   6688: out<=1;
   6689: out<=1;
   6690: out<=1;
   6691: out<=1;
   6692: out<=0;
   6693: out<=1;
   6694: out<=1;
   6695: out<=0;
   6696: out<=0;
   6697: out<=1;
   6698: out<=0;
   6699: out<=1;
   6700: out<=1;
   6701: out<=1;
   6702: out<=0;
   6703: out<=0;
   6704: out<=1;
   6705: out<=0;
   6706: out<=0;
   6707: out<=1;
   6708: out<=1;
   6709: out<=1;
   6710: out<=1;
   6711: out<=1;
   6712: out<=1;
   6713: out<=1;
   6714: out<=0;
   6715: out<=0;
   6716: out<=1;
   6717: out<=0;
   6718: out<=1;
   6719: out<=0;
   6720: out<=0;
   6721: out<=1;
   6722: out<=0;
   6723: out<=1;
   6724: out<=0;
   6725: out<=0;
   6726: out<=1;
   6727: out<=1;
   6728: out<=1;
   6729: out<=1;
   6730: out<=1;
   6731: out<=1;
   6732: out<=1;
   6733: out<=0;
   6734: out<=0;
   6735: out<=1;
   6736: out<=1;
   6737: out<=1;
   6738: out<=0;
   6739: out<=0;
   6740: out<=0;
   6741: out<=1;
   6742: out<=0;
   6743: out<=1;
   6744: out<=1;
   6745: out<=0;
   6746: out<=0;
   6747: out<=1;
   6748: out<=0;
   6749: out<=0;
   6750: out<=0;
   6751: out<=0;
   6752: out<=1;
   6753: out<=1;
   6754: out<=1;
   6755: out<=1;
   6756: out<=0;
   6757: out<=1;
   6758: out<=1;
   6759: out<=0;
   6760: out<=0;
   6761: out<=1;
   6762: out<=0;
   6763: out<=1;
   6764: out<=1;
   6765: out<=1;
   6766: out<=0;
   6767: out<=0;
   6768: out<=0;
   6769: out<=1;
   6770: out<=1;
   6771: out<=0;
   6772: out<=0;
   6773: out<=0;
   6774: out<=0;
   6775: out<=0;
   6776: out<=0;
   6777: out<=0;
   6778: out<=1;
   6779: out<=1;
   6780: out<=0;
   6781: out<=1;
   6782: out<=0;
   6783: out<=1;
   6784: out<=1;
   6785: out<=0;
   6786: out<=1;
   6787: out<=0;
   6788: out<=1;
   6789: out<=1;
   6790: out<=0;
   6791: out<=0;
   6792: out<=0;
   6793: out<=0;
   6794: out<=0;
   6795: out<=0;
   6796: out<=0;
   6797: out<=1;
   6798: out<=1;
   6799: out<=0;
   6800: out<=0;
   6801: out<=0;
   6802: out<=1;
   6803: out<=1;
   6804: out<=1;
   6805: out<=0;
   6806: out<=1;
   6807: out<=0;
   6808: out<=0;
   6809: out<=1;
   6810: out<=1;
   6811: out<=0;
   6812: out<=1;
   6813: out<=1;
   6814: out<=1;
   6815: out<=1;
   6816: out<=1;
   6817: out<=1;
   6818: out<=1;
   6819: out<=1;
   6820: out<=0;
   6821: out<=1;
   6822: out<=1;
   6823: out<=0;
   6824: out<=0;
   6825: out<=1;
   6826: out<=0;
   6827: out<=1;
   6828: out<=1;
   6829: out<=1;
   6830: out<=0;
   6831: out<=0;
   6832: out<=0;
   6833: out<=1;
   6834: out<=1;
   6835: out<=0;
   6836: out<=0;
   6837: out<=0;
   6838: out<=0;
   6839: out<=0;
   6840: out<=0;
   6841: out<=0;
   6842: out<=1;
   6843: out<=1;
   6844: out<=0;
   6845: out<=1;
   6846: out<=0;
   6847: out<=1;
   6848: out<=0;
   6849: out<=1;
   6850: out<=0;
   6851: out<=1;
   6852: out<=0;
   6853: out<=0;
   6854: out<=1;
   6855: out<=1;
   6856: out<=1;
   6857: out<=1;
   6858: out<=1;
   6859: out<=1;
   6860: out<=1;
   6861: out<=0;
   6862: out<=0;
   6863: out<=1;
   6864: out<=0;
   6865: out<=0;
   6866: out<=1;
   6867: out<=1;
   6868: out<=1;
   6869: out<=0;
   6870: out<=1;
   6871: out<=0;
   6872: out<=0;
   6873: out<=1;
   6874: out<=1;
   6875: out<=0;
   6876: out<=1;
   6877: out<=1;
   6878: out<=1;
   6879: out<=1;
   6880: out<=1;
   6881: out<=1;
   6882: out<=1;
   6883: out<=1;
   6884: out<=0;
   6885: out<=1;
   6886: out<=1;
   6887: out<=0;
   6888: out<=0;
   6889: out<=1;
   6890: out<=0;
   6891: out<=1;
   6892: out<=1;
   6893: out<=1;
   6894: out<=0;
   6895: out<=0;
   6896: out<=1;
   6897: out<=0;
   6898: out<=0;
   6899: out<=1;
   6900: out<=1;
   6901: out<=1;
   6902: out<=1;
   6903: out<=1;
   6904: out<=1;
   6905: out<=1;
   6906: out<=0;
   6907: out<=0;
   6908: out<=1;
   6909: out<=0;
   6910: out<=1;
   6911: out<=0;
   6912: out<=1;
   6913: out<=1;
   6914: out<=0;
   6915: out<=0;
   6916: out<=0;
   6917: out<=1;
   6918: out<=0;
   6919: out<=1;
   6920: out<=1;
   6921: out<=0;
   6922: out<=0;
   6923: out<=1;
   6924: out<=0;
   6925: out<=0;
   6926: out<=0;
   6927: out<=0;
   6928: out<=0;
   6929: out<=1;
   6930: out<=0;
   6931: out<=1;
   6932: out<=0;
   6933: out<=0;
   6934: out<=1;
   6935: out<=1;
   6936: out<=1;
   6937: out<=1;
   6938: out<=1;
   6939: out<=1;
   6940: out<=1;
   6941: out<=0;
   6942: out<=0;
   6943: out<=1;
   6944: out<=0;
   6945: out<=1;
   6946: out<=1;
   6947: out<=0;
   6948: out<=0;
   6949: out<=0;
   6950: out<=0;
   6951: out<=0;
   6952: out<=0;
   6953: out<=0;
   6954: out<=1;
   6955: out<=1;
   6956: out<=0;
   6957: out<=1;
   6958: out<=0;
   6959: out<=1;
   6960: out<=1;
   6961: out<=1;
   6962: out<=1;
   6963: out<=1;
   6964: out<=0;
   6965: out<=1;
   6966: out<=1;
   6967: out<=0;
   6968: out<=0;
   6969: out<=1;
   6970: out<=0;
   6971: out<=1;
   6972: out<=1;
   6973: out<=1;
   6974: out<=0;
   6975: out<=0;
   6976: out<=1;
   6977: out<=1;
   6978: out<=0;
   6979: out<=0;
   6980: out<=0;
   6981: out<=1;
   6982: out<=0;
   6983: out<=1;
   6984: out<=1;
   6985: out<=0;
   6986: out<=0;
   6987: out<=1;
   6988: out<=0;
   6989: out<=0;
   6990: out<=0;
   6991: out<=0;
   6992: out<=1;
   6993: out<=0;
   6994: out<=1;
   6995: out<=0;
   6996: out<=1;
   6997: out<=1;
   6998: out<=0;
   6999: out<=0;
   7000: out<=0;
   7001: out<=0;
   7002: out<=0;
   7003: out<=0;
   7004: out<=0;
   7005: out<=1;
   7006: out<=1;
   7007: out<=0;
   7008: out<=1;
   7009: out<=0;
   7010: out<=0;
   7011: out<=1;
   7012: out<=1;
   7013: out<=1;
   7014: out<=1;
   7015: out<=1;
   7016: out<=1;
   7017: out<=1;
   7018: out<=0;
   7019: out<=0;
   7020: out<=1;
   7021: out<=0;
   7022: out<=1;
   7023: out<=0;
   7024: out<=1;
   7025: out<=1;
   7026: out<=1;
   7027: out<=1;
   7028: out<=0;
   7029: out<=1;
   7030: out<=1;
   7031: out<=0;
   7032: out<=0;
   7033: out<=1;
   7034: out<=0;
   7035: out<=1;
   7036: out<=1;
   7037: out<=1;
   7038: out<=0;
   7039: out<=0;
   7040: out<=0;
   7041: out<=0;
   7042: out<=1;
   7043: out<=1;
   7044: out<=1;
   7045: out<=0;
   7046: out<=1;
   7047: out<=0;
   7048: out<=0;
   7049: out<=1;
   7050: out<=1;
   7051: out<=0;
   7052: out<=1;
   7053: out<=1;
   7054: out<=1;
   7055: out<=1;
   7056: out<=0;
   7057: out<=1;
   7058: out<=0;
   7059: out<=1;
   7060: out<=0;
   7061: out<=0;
   7062: out<=1;
   7063: out<=1;
   7064: out<=1;
   7065: out<=1;
   7066: out<=1;
   7067: out<=1;
   7068: out<=1;
   7069: out<=0;
   7070: out<=0;
   7071: out<=1;
   7072: out<=1;
   7073: out<=0;
   7074: out<=0;
   7075: out<=1;
   7076: out<=1;
   7077: out<=1;
   7078: out<=1;
   7079: out<=1;
   7080: out<=1;
   7081: out<=1;
   7082: out<=0;
   7083: out<=0;
   7084: out<=1;
   7085: out<=0;
   7086: out<=1;
   7087: out<=0;
   7088: out<=1;
   7089: out<=1;
   7090: out<=1;
   7091: out<=1;
   7092: out<=0;
   7093: out<=1;
   7094: out<=1;
   7095: out<=0;
   7096: out<=0;
   7097: out<=1;
   7098: out<=0;
   7099: out<=1;
   7100: out<=1;
   7101: out<=1;
   7102: out<=0;
   7103: out<=0;
   7104: out<=0;
   7105: out<=0;
   7106: out<=1;
   7107: out<=1;
   7108: out<=1;
   7109: out<=0;
   7110: out<=1;
   7111: out<=0;
   7112: out<=0;
   7113: out<=1;
   7114: out<=1;
   7115: out<=0;
   7116: out<=1;
   7117: out<=1;
   7118: out<=1;
   7119: out<=1;
   7120: out<=1;
   7121: out<=0;
   7122: out<=1;
   7123: out<=0;
   7124: out<=1;
   7125: out<=1;
   7126: out<=0;
   7127: out<=0;
   7128: out<=0;
   7129: out<=0;
   7130: out<=0;
   7131: out<=0;
   7132: out<=0;
   7133: out<=1;
   7134: out<=1;
   7135: out<=0;
   7136: out<=0;
   7137: out<=1;
   7138: out<=1;
   7139: out<=0;
   7140: out<=0;
   7141: out<=0;
   7142: out<=0;
   7143: out<=0;
   7144: out<=0;
   7145: out<=0;
   7146: out<=1;
   7147: out<=1;
   7148: out<=0;
   7149: out<=1;
   7150: out<=0;
   7151: out<=1;
   7152: out<=1;
   7153: out<=1;
   7154: out<=1;
   7155: out<=1;
   7156: out<=0;
   7157: out<=1;
   7158: out<=1;
   7159: out<=0;
   7160: out<=0;
   7161: out<=1;
   7162: out<=0;
   7163: out<=1;
   7164: out<=1;
   7165: out<=1;
   7166: out<=0;
   7167: out<=0;
   7168: out<=0;
   7169: out<=1;
   7170: out<=1;
   7171: out<=0;
   7172: out<=1;
   7173: out<=1;
   7174: out<=1;
   7175: out<=1;
   7176: out<=1;
   7177: out<=1;
   7178: out<=0;
   7179: out<=0;
   7180: out<=0;
   7181: out<=1;
   7182: out<=0;
   7183: out<=1;
   7184: out<=1;
   7185: out<=1;
   7186: out<=1;
   7187: out<=1;
   7188: out<=1;
   7189: out<=0;
   7190: out<=0;
   7191: out<=1;
   7192: out<=1;
   7193: out<=0;
   7194: out<=1;
   7195: out<=0;
   7196: out<=1;
   7197: out<=1;
   7198: out<=0;
   7199: out<=0;
   7200: out<=0;
   7201: out<=0;
   7202: out<=1;
   7203: out<=1;
   7204: out<=0;
   7205: out<=1;
   7206: out<=0;
   7207: out<=1;
   7208: out<=1;
   7209: out<=0;
   7210: out<=0;
   7211: out<=1;
   7212: out<=1;
   7213: out<=1;
   7214: out<=1;
   7215: out<=1;
   7216: out<=1;
   7217: out<=0;
   7218: out<=1;
   7219: out<=0;
   7220: out<=0;
   7221: out<=0;
   7222: out<=1;
   7223: out<=1;
   7224: out<=1;
   7225: out<=1;
   7226: out<=1;
   7227: out<=1;
   7228: out<=0;
   7229: out<=1;
   7230: out<=1;
   7231: out<=0;
   7232: out<=1;
   7233: out<=0;
   7234: out<=0;
   7235: out<=1;
   7236: out<=0;
   7237: out<=0;
   7238: out<=0;
   7239: out<=0;
   7240: out<=0;
   7241: out<=0;
   7242: out<=1;
   7243: out<=1;
   7244: out<=1;
   7245: out<=0;
   7246: out<=1;
   7247: out<=0;
   7248: out<=1;
   7249: out<=1;
   7250: out<=1;
   7251: out<=1;
   7252: out<=1;
   7253: out<=0;
   7254: out<=0;
   7255: out<=1;
   7256: out<=1;
   7257: out<=0;
   7258: out<=1;
   7259: out<=0;
   7260: out<=1;
   7261: out<=1;
   7262: out<=0;
   7263: out<=0;
   7264: out<=0;
   7265: out<=0;
   7266: out<=1;
   7267: out<=1;
   7268: out<=0;
   7269: out<=1;
   7270: out<=0;
   7271: out<=1;
   7272: out<=1;
   7273: out<=0;
   7274: out<=0;
   7275: out<=1;
   7276: out<=1;
   7277: out<=1;
   7278: out<=1;
   7279: out<=1;
   7280: out<=0;
   7281: out<=1;
   7282: out<=0;
   7283: out<=1;
   7284: out<=1;
   7285: out<=1;
   7286: out<=0;
   7287: out<=0;
   7288: out<=0;
   7289: out<=0;
   7290: out<=0;
   7291: out<=0;
   7292: out<=1;
   7293: out<=0;
   7294: out<=0;
   7295: out<=1;
   7296: out<=1;
   7297: out<=0;
   7298: out<=0;
   7299: out<=1;
   7300: out<=0;
   7301: out<=0;
   7302: out<=0;
   7303: out<=0;
   7304: out<=0;
   7305: out<=0;
   7306: out<=1;
   7307: out<=1;
   7308: out<=1;
   7309: out<=0;
   7310: out<=1;
   7311: out<=0;
   7312: out<=1;
   7313: out<=1;
   7314: out<=1;
   7315: out<=1;
   7316: out<=1;
   7317: out<=0;
   7318: out<=0;
   7319: out<=1;
   7320: out<=1;
   7321: out<=0;
   7322: out<=1;
   7323: out<=0;
   7324: out<=1;
   7325: out<=1;
   7326: out<=0;
   7327: out<=0;
   7328: out<=1;
   7329: out<=1;
   7330: out<=0;
   7331: out<=0;
   7332: out<=1;
   7333: out<=0;
   7334: out<=1;
   7335: out<=0;
   7336: out<=0;
   7337: out<=1;
   7338: out<=1;
   7339: out<=0;
   7340: out<=0;
   7341: out<=0;
   7342: out<=0;
   7343: out<=0;
   7344: out<=1;
   7345: out<=0;
   7346: out<=1;
   7347: out<=0;
   7348: out<=0;
   7349: out<=0;
   7350: out<=1;
   7351: out<=1;
   7352: out<=1;
   7353: out<=1;
   7354: out<=1;
   7355: out<=1;
   7356: out<=0;
   7357: out<=1;
   7358: out<=1;
   7359: out<=0;
   7360: out<=0;
   7361: out<=1;
   7362: out<=1;
   7363: out<=0;
   7364: out<=1;
   7365: out<=1;
   7366: out<=1;
   7367: out<=1;
   7368: out<=1;
   7369: out<=1;
   7370: out<=0;
   7371: out<=0;
   7372: out<=0;
   7373: out<=1;
   7374: out<=0;
   7375: out<=1;
   7376: out<=1;
   7377: out<=1;
   7378: out<=1;
   7379: out<=1;
   7380: out<=1;
   7381: out<=0;
   7382: out<=0;
   7383: out<=1;
   7384: out<=1;
   7385: out<=0;
   7386: out<=1;
   7387: out<=0;
   7388: out<=1;
   7389: out<=1;
   7390: out<=0;
   7391: out<=0;
   7392: out<=1;
   7393: out<=1;
   7394: out<=0;
   7395: out<=0;
   7396: out<=1;
   7397: out<=0;
   7398: out<=1;
   7399: out<=0;
   7400: out<=0;
   7401: out<=1;
   7402: out<=1;
   7403: out<=0;
   7404: out<=0;
   7405: out<=0;
   7406: out<=0;
   7407: out<=0;
   7408: out<=0;
   7409: out<=1;
   7410: out<=0;
   7411: out<=1;
   7412: out<=1;
   7413: out<=1;
   7414: out<=0;
   7415: out<=0;
   7416: out<=0;
   7417: out<=0;
   7418: out<=0;
   7419: out<=0;
   7420: out<=1;
   7421: out<=0;
   7422: out<=0;
   7423: out<=1;
   7424: out<=1;
   7425: out<=1;
   7426: out<=1;
   7427: out<=1;
   7428: out<=1;
   7429: out<=0;
   7430: out<=0;
   7431: out<=1;
   7432: out<=1;
   7433: out<=0;
   7434: out<=1;
   7435: out<=0;
   7436: out<=1;
   7437: out<=1;
   7438: out<=0;
   7439: out<=0;
   7440: out<=1;
   7441: out<=0;
   7442: out<=0;
   7443: out<=1;
   7444: out<=0;
   7445: out<=0;
   7446: out<=0;
   7447: out<=0;
   7448: out<=0;
   7449: out<=0;
   7450: out<=1;
   7451: out<=1;
   7452: out<=1;
   7453: out<=0;
   7454: out<=1;
   7455: out<=0;
   7456: out<=0;
   7457: out<=1;
   7458: out<=0;
   7459: out<=1;
   7460: out<=1;
   7461: out<=1;
   7462: out<=0;
   7463: out<=0;
   7464: out<=0;
   7465: out<=0;
   7466: out<=0;
   7467: out<=0;
   7468: out<=1;
   7469: out<=0;
   7470: out<=0;
   7471: out<=1;
   7472: out<=0;
   7473: out<=0;
   7474: out<=1;
   7475: out<=1;
   7476: out<=0;
   7477: out<=1;
   7478: out<=0;
   7479: out<=1;
   7480: out<=1;
   7481: out<=0;
   7482: out<=0;
   7483: out<=1;
   7484: out<=1;
   7485: out<=1;
   7486: out<=1;
   7487: out<=1;
   7488: out<=1;
   7489: out<=1;
   7490: out<=1;
   7491: out<=1;
   7492: out<=1;
   7493: out<=0;
   7494: out<=0;
   7495: out<=1;
   7496: out<=1;
   7497: out<=0;
   7498: out<=1;
   7499: out<=0;
   7500: out<=1;
   7501: out<=1;
   7502: out<=0;
   7503: out<=0;
   7504: out<=0;
   7505: out<=1;
   7506: out<=1;
   7507: out<=0;
   7508: out<=1;
   7509: out<=1;
   7510: out<=1;
   7511: out<=1;
   7512: out<=1;
   7513: out<=1;
   7514: out<=0;
   7515: out<=0;
   7516: out<=0;
   7517: out<=1;
   7518: out<=0;
   7519: out<=1;
   7520: out<=1;
   7521: out<=0;
   7522: out<=1;
   7523: out<=0;
   7524: out<=0;
   7525: out<=0;
   7526: out<=1;
   7527: out<=1;
   7528: out<=1;
   7529: out<=1;
   7530: out<=1;
   7531: out<=1;
   7532: out<=0;
   7533: out<=1;
   7534: out<=1;
   7535: out<=0;
   7536: out<=0;
   7537: out<=0;
   7538: out<=1;
   7539: out<=1;
   7540: out<=0;
   7541: out<=1;
   7542: out<=0;
   7543: out<=1;
   7544: out<=1;
   7545: out<=0;
   7546: out<=0;
   7547: out<=1;
   7548: out<=1;
   7549: out<=1;
   7550: out<=1;
   7551: out<=1;
   7552: out<=1;
   7553: out<=1;
   7554: out<=1;
   7555: out<=1;
   7556: out<=1;
   7557: out<=0;
   7558: out<=0;
   7559: out<=1;
   7560: out<=1;
   7561: out<=0;
   7562: out<=1;
   7563: out<=0;
   7564: out<=1;
   7565: out<=1;
   7566: out<=0;
   7567: out<=0;
   7568: out<=0;
   7569: out<=1;
   7570: out<=1;
   7571: out<=0;
   7572: out<=1;
   7573: out<=1;
   7574: out<=1;
   7575: out<=1;
   7576: out<=1;
   7577: out<=1;
   7578: out<=0;
   7579: out<=0;
   7580: out<=0;
   7581: out<=1;
   7582: out<=0;
   7583: out<=1;
   7584: out<=0;
   7585: out<=1;
   7586: out<=0;
   7587: out<=1;
   7588: out<=1;
   7589: out<=1;
   7590: out<=0;
   7591: out<=0;
   7592: out<=0;
   7593: out<=0;
   7594: out<=0;
   7595: out<=0;
   7596: out<=1;
   7597: out<=0;
   7598: out<=0;
   7599: out<=1;
   7600: out<=1;
   7601: out<=1;
   7602: out<=0;
   7603: out<=0;
   7604: out<=1;
   7605: out<=0;
   7606: out<=1;
   7607: out<=0;
   7608: out<=0;
   7609: out<=1;
   7610: out<=1;
   7611: out<=0;
   7612: out<=0;
   7613: out<=0;
   7614: out<=0;
   7615: out<=0;
   7616: out<=1;
   7617: out<=1;
   7618: out<=1;
   7619: out<=1;
   7620: out<=1;
   7621: out<=0;
   7622: out<=0;
   7623: out<=1;
   7624: out<=1;
   7625: out<=0;
   7626: out<=1;
   7627: out<=0;
   7628: out<=1;
   7629: out<=1;
   7630: out<=0;
   7631: out<=0;
   7632: out<=1;
   7633: out<=0;
   7634: out<=0;
   7635: out<=1;
   7636: out<=0;
   7637: out<=0;
   7638: out<=0;
   7639: out<=0;
   7640: out<=0;
   7641: out<=0;
   7642: out<=1;
   7643: out<=1;
   7644: out<=1;
   7645: out<=0;
   7646: out<=1;
   7647: out<=0;
   7648: out<=1;
   7649: out<=0;
   7650: out<=1;
   7651: out<=0;
   7652: out<=0;
   7653: out<=0;
   7654: out<=1;
   7655: out<=1;
   7656: out<=1;
   7657: out<=1;
   7658: out<=1;
   7659: out<=1;
   7660: out<=0;
   7661: out<=1;
   7662: out<=1;
   7663: out<=0;
   7664: out<=1;
   7665: out<=1;
   7666: out<=0;
   7667: out<=0;
   7668: out<=1;
   7669: out<=0;
   7670: out<=1;
   7671: out<=0;
   7672: out<=0;
   7673: out<=1;
   7674: out<=1;
   7675: out<=0;
   7676: out<=0;
   7677: out<=0;
   7678: out<=0;
   7679: out<=0;
   7680: out<=1;
   7681: out<=1;
   7682: out<=0;
   7683: out<=0;
   7684: out<=1;
   7685: out<=0;
   7686: out<=1;
   7687: out<=0;
   7688: out<=0;
   7689: out<=1;
   7690: out<=1;
   7691: out<=0;
   7692: out<=0;
   7693: out<=0;
   7694: out<=0;
   7695: out<=0;
   7696: out<=1;
   7697: out<=0;
   7698: out<=1;
   7699: out<=0;
   7700: out<=0;
   7701: out<=0;
   7702: out<=1;
   7703: out<=1;
   7704: out<=1;
   7705: out<=1;
   7706: out<=1;
   7707: out<=1;
   7708: out<=0;
   7709: out<=1;
   7710: out<=1;
   7711: out<=0;
   7712: out<=1;
   7713: out<=0;
   7714: out<=0;
   7715: out<=1;
   7716: out<=0;
   7717: out<=0;
   7718: out<=0;
   7719: out<=0;
   7720: out<=0;
   7721: out<=0;
   7722: out<=1;
   7723: out<=1;
   7724: out<=1;
   7725: out<=0;
   7726: out<=1;
   7727: out<=0;
   7728: out<=1;
   7729: out<=1;
   7730: out<=1;
   7731: out<=1;
   7732: out<=1;
   7733: out<=0;
   7734: out<=0;
   7735: out<=1;
   7736: out<=1;
   7737: out<=0;
   7738: out<=1;
   7739: out<=0;
   7740: out<=1;
   7741: out<=1;
   7742: out<=0;
   7743: out<=0;
   7744: out<=1;
   7745: out<=1;
   7746: out<=0;
   7747: out<=0;
   7748: out<=1;
   7749: out<=0;
   7750: out<=1;
   7751: out<=0;
   7752: out<=0;
   7753: out<=1;
   7754: out<=1;
   7755: out<=0;
   7756: out<=0;
   7757: out<=0;
   7758: out<=0;
   7759: out<=0;
   7760: out<=0;
   7761: out<=1;
   7762: out<=0;
   7763: out<=1;
   7764: out<=1;
   7765: out<=1;
   7766: out<=0;
   7767: out<=0;
   7768: out<=0;
   7769: out<=0;
   7770: out<=0;
   7771: out<=0;
   7772: out<=1;
   7773: out<=0;
   7774: out<=0;
   7775: out<=1;
   7776: out<=0;
   7777: out<=1;
   7778: out<=1;
   7779: out<=0;
   7780: out<=1;
   7781: out<=1;
   7782: out<=1;
   7783: out<=1;
   7784: out<=1;
   7785: out<=1;
   7786: out<=0;
   7787: out<=0;
   7788: out<=0;
   7789: out<=1;
   7790: out<=0;
   7791: out<=1;
   7792: out<=1;
   7793: out<=1;
   7794: out<=1;
   7795: out<=1;
   7796: out<=1;
   7797: out<=0;
   7798: out<=0;
   7799: out<=1;
   7800: out<=1;
   7801: out<=0;
   7802: out<=1;
   7803: out<=0;
   7804: out<=1;
   7805: out<=1;
   7806: out<=0;
   7807: out<=0;
   7808: out<=0;
   7809: out<=0;
   7810: out<=1;
   7811: out<=1;
   7812: out<=0;
   7813: out<=1;
   7814: out<=0;
   7815: out<=1;
   7816: out<=1;
   7817: out<=0;
   7818: out<=0;
   7819: out<=1;
   7820: out<=1;
   7821: out<=1;
   7822: out<=1;
   7823: out<=1;
   7824: out<=1;
   7825: out<=0;
   7826: out<=1;
   7827: out<=0;
   7828: out<=0;
   7829: out<=0;
   7830: out<=1;
   7831: out<=1;
   7832: out<=1;
   7833: out<=1;
   7834: out<=1;
   7835: out<=1;
   7836: out<=0;
   7837: out<=1;
   7838: out<=1;
   7839: out<=0;
   7840: out<=0;
   7841: out<=1;
   7842: out<=1;
   7843: out<=0;
   7844: out<=1;
   7845: out<=1;
   7846: out<=1;
   7847: out<=1;
   7848: out<=1;
   7849: out<=1;
   7850: out<=0;
   7851: out<=0;
   7852: out<=0;
   7853: out<=1;
   7854: out<=0;
   7855: out<=1;
   7856: out<=1;
   7857: out<=1;
   7858: out<=1;
   7859: out<=1;
   7860: out<=1;
   7861: out<=0;
   7862: out<=0;
   7863: out<=1;
   7864: out<=1;
   7865: out<=0;
   7866: out<=1;
   7867: out<=0;
   7868: out<=1;
   7869: out<=1;
   7870: out<=0;
   7871: out<=0;
   7872: out<=0;
   7873: out<=0;
   7874: out<=1;
   7875: out<=1;
   7876: out<=0;
   7877: out<=1;
   7878: out<=0;
   7879: out<=1;
   7880: out<=1;
   7881: out<=0;
   7882: out<=0;
   7883: out<=1;
   7884: out<=1;
   7885: out<=1;
   7886: out<=1;
   7887: out<=1;
   7888: out<=0;
   7889: out<=1;
   7890: out<=0;
   7891: out<=1;
   7892: out<=1;
   7893: out<=1;
   7894: out<=0;
   7895: out<=0;
   7896: out<=0;
   7897: out<=0;
   7898: out<=0;
   7899: out<=0;
   7900: out<=1;
   7901: out<=0;
   7902: out<=0;
   7903: out<=1;
   7904: out<=1;
   7905: out<=0;
   7906: out<=0;
   7907: out<=1;
   7908: out<=0;
   7909: out<=0;
   7910: out<=0;
   7911: out<=0;
   7912: out<=0;
   7913: out<=0;
   7914: out<=1;
   7915: out<=1;
   7916: out<=1;
   7917: out<=0;
   7918: out<=1;
   7919: out<=0;
   7920: out<=1;
   7921: out<=1;
   7922: out<=1;
   7923: out<=1;
   7924: out<=1;
   7925: out<=0;
   7926: out<=0;
   7927: out<=1;
   7928: out<=1;
   7929: out<=0;
   7930: out<=1;
   7931: out<=0;
   7932: out<=1;
   7933: out<=1;
   7934: out<=0;
   7935: out<=0;
   7936: out<=0;
   7937: out<=1;
   7938: out<=0;
   7939: out<=1;
   7940: out<=1;
   7941: out<=1;
   7942: out<=0;
   7943: out<=0;
   7944: out<=0;
   7945: out<=0;
   7946: out<=0;
   7947: out<=0;
   7948: out<=1;
   7949: out<=0;
   7950: out<=0;
   7951: out<=1;
   7952: out<=1;
   7953: out<=1;
   7954: out<=0;
   7955: out<=0;
   7956: out<=1;
   7957: out<=0;
   7958: out<=1;
   7959: out<=0;
   7960: out<=0;
   7961: out<=1;
   7962: out<=1;
   7963: out<=0;
   7964: out<=0;
   7965: out<=0;
   7966: out<=0;
   7967: out<=0;
   7968: out<=1;
   7969: out<=1;
   7970: out<=1;
   7971: out<=1;
   7972: out<=1;
   7973: out<=0;
   7974: out<=0;
   7975: out<=1;
   7976: out<=1;
   7977: out<=0;
   7978: out<=1;
   7979: out<=0;
   7980: out<=1;
   7981: out<=1;
   7982: out<=0;
   7983: out<=0;
   7984: out<=0;
   7985: out<=1;
   7986: out<=1;
   7987: out<=0;
   7988: out<=1;
   7989: out<=1;
   7990: out<=1;
   7991: out<=1;
   7992: out<=1;
   7993: out<=1;
   7994: out<=0;
   7995: out<=0;
   7996: out<=0;
   7997: out<=1;
   7998: out<=0;
   7999: out<=1;
   8000: out<=1;
   8001: out<=0;
   8002: out<=1;
   8003: out<=0;
   8004: out<=0;
   8005: out<=0;
   8006: out<=1;
   8007: out<=1;
   8008: out<=1;
   8009: out<=1;
   8010: out<=1;
   8011: out<=1;
   8012: out<=0;
   8013: out<=1;
   8014: out<=1;
   8015: out<=0;
   8016: out<=1;
   8017: out<=1;
   8018: out<=0;
   8019: out<=0;
   8020: out<=1;
   8021: out<=0;
   8022: out<=1;
   8023: out<=0;
   8024: out<=0;
   8025: out<=1;
   8026: out<=1;
   8027: out<=0;
   8028: out<=0;
   8029: out<=0;
   8030: out<=0;
   8031: out<=0;
   8032: out<=1;
   8033: out<=1;
   8034: out<=1;
   8035: out<=1;
   8036: out<=1;
   8037: out<=0;
   8038: out<=0;
   8039: out<=1;
   8040: out<=1;
   8041: out<=0;
   8042: out<=1;
   8043: out<=0;
   8044: out<=1;
   8045: out<=1;
   8046: out<=0;
   8047: out<=0;
   8048: out<=1;
   8049: out<=0;
   8050: out<=0;
   8051: out<=1;
   8052: out<=0;
   8053: out<=0;
   8054: out<=0;
   8055: out<=0;
   8056: out<=0;
   8057: out<=0;
   8058: out<=1;
   8059: out<=1;
   8060: out<=1;
   8061: out<=0;
   8062: out<=1;
   8063: out<=0;
   8064: out<=0;
   8065: out<=1;
   8066: out<=0;
   8067: out<=1;
   8068: out<=1;
   8069: out<=1;
   8070: out<=0;
   8071: out<=0;
   8072: out<=0;
   8073: out<=0;
   8074: out<=0;
   8075: out<=0;
   8076: out<=1;
   8077: out<=0;
   8078: out<=0;
   8079: out<=1;
   8080: out<=0;
   8081: out<=0;
   8082: out<=1;
   8083: out<=1;
   8084: out<=0;
   8085: out<=1;
   8086: out<=0;
   8087: out<=1;
   8088: out<=1;
   8089: out<=0;
   8090: out<=0;
   8091: out<=1;
   8092: out<=1;
   8093: out<=1;
   8094: out<=1;
   8095: out<=1;
   8096: out<=1;
   8097: out<=1;
   8098: out<=1;
   8099: out<=1;
   8100: out<=1;
   8101: out<=0;
   8102: out<=0;
   8103: out<=1;
   8104: out<=1;
   8105: out<=0;
   8106: out<=1;
   8107: out<=0;
   8108: out<=1;
   8109: out<=1;
   8110: out<=0;
   8111: out<=0;
   8112: out<=1;
   8113: out<=0;
   8114: out<=0;
   8115: out<=1;
   8116: out<=0;
   8117: out<=0;
   8118: out<=0;
   8119: out<=0;
   8120: out<=0;
   8121: out<=0;
   8122: out<=1;
   8123: out<=1;
   8124: out<=1;
   8125: out<=0;
   8126: out<=1;
   8127: out<=0;
   8128: out<=1;
   8129: out<=0;
   8130: out<=1;
   8131: out<=0;
   8132: out<=0;
   8133: out<=0;
   8134: out<=1;
   8135: out<=1;
   8136: out<=1;
   8137: out<=1;
   8138: out<=1;
   8139: out<=1;
   8140: out<=0;
   8141: out<=1;
   8142: out<=1;
   8143: out<=0;
   8144: out<=0;
   8145: out<=0;
   8146: out<=1;
   8147: out<=1;
   8148: out<=0;
   8149: out<=1;
   8150: out<=0;
   8151: out<=1;
   8152: out<=1;
   8153: out<=0;
   8154: out<=0;
   8155: out<=1;
   8156: out<=1;
   8157: out<=1;
   8158: out<=1;
   8159: out<=1;
   8160: out<=1;
   8161: out<=1;
   8162: out<=1;
   8163: out<=1;
   8164: out<=1;
   8165: out<=0;
   8166: out<=0;
   8167: out<=1;
   8168: out<=1;
   8169: out<=0;
   8170: out<=1;
   8171: out<=0;
   8172: out<=1;
   8173: out<=1;
   8174: out<=0;
   8175: out<=0;
   8176: out<=0;
   8177: out<=1;
   8178: out<=1;
   8179: out<=0;
   8180: out<=1;
   8181: out<=1;
   8182: out<=1;
   8183: out<=1;
   8184: out<=1;
   8185: out<=1;
   8186: out<=0;
   8187: out<=0;
   8188: out<=0;
   8189: out<=1;
   8190: out<=0;
   8191: out<=1;
   8192: out<=0;
   8193: out<=1;
   8194: out<=0;
   8195: out<=1;
   8196: out<=1;
   8197: out<=1;
   8198: out<=0;
   8199: out<=0;
   8200: out<=0;
   8201: out<=0;
   8202: out<=0;
   8203: out<=0;
   8204: out<=1;
   8205: out<=0;
   8206: out<=0;
   8207: out<=1;
   8208: out<=1;
   8209: out<=1;
   8210: out<=0;
   8211: out<=0;
   8212: out<=1;
   8213: out<=0;
   8214: out<=1;
   8215: out<=0;
   8216: out<=0;
   8217: out<=1;
   8218: out<=1;
   8219: out<=0;
   8220: out<=0;
   8221: out<=0;
   8222: out<=0;
   8223: out<=0;
   8224: out<=0;
   8225: out<=0;
   8226: out<=0;
   8227: out<=0;
   8228: out<=0;
   8229: out<=1;
   8230: out<=1;
   8231: out<=0;
   8232: out<=0;
   8233: out<=1;
   8234: out<=0;
   8235: out<=1;
   8236: out<=0;
   8237: out<=0;
   8238: out<=1;
   8239: out<=1;
   8240: out<=1;
   8241: out<=0;
   8242: out<=0;
   8243: out<=1;
   8244: out<=0;
   8245: out<=0;
   8246: out<=0;
   8247: out<=0;
   8248: out<=0;
   8249: out<=0;
   8250: out<=1;
   8251: out<=1;
   8252: out<=1;
   8253: out<=0;
   8254: out<=1;
   8255: out<=0;
   8256: out<=1;
   8257: out<=0;
   8258: out<=1;
   8259: out<=0;
   8260: out<=0;
   8261: out<=0;
   8262: out<=1;
   8263: out<=1;
   8264: out<=1;
   8265: out<=1;
   8266: out<=1;
   8267: out<=1;
   8268: out<=0;
   8269: out<=1;
   8270: out<=1;
   8271: out<=0;
   8272: out<=1;
   8273: out<=1;
   8274: out<=0;
   8275: out<=0;
   8276: out<=1;
   8277: out<=0;
   8278: out<=1;
   8279: out<=0;
   8280: out<=0;
   8281: out<=1;
   8282: out<=1;
   8283: out<=0;
   8284: out<=0;
   8285: out<=0;
   8286: out<=0;
   8287: out<=0;
   8288: out<=0;
   8289: out<=0;
   8290: out<=0;
   8291: out<=0;
   8292: out<=0;
   8293: out<=1;
   8294: out<=1;
   8295: out<=0;
   8296: out<=0;
   8297: out<=1;
   8298: out<=0;
   8299: out<=1;
   8300: out<=0;
   8301: out<=0;
   8302: out<=1;
   8303: out<=1;
   8304: out<=0;
   8305: out<=1;
   8306: out<=1;
   8307: out<=0;
   8308: out<=1;
   8309: out<=1;
   8310: out<=1;
   8311: out<=1;
   8312: out<=1;
   8313: out<=1;
   8314: out<=0;
   8315: out<=0;
   8316: out<=0;
   8317: out<=1;
   8318: out<=0;
   8319: out<=1;
   8320: out<=0;
   8321: out<=1;
   8322: out<=0;
   8323: out<=1;
   8324: out<=1;
   8325: out<=1;
   8326: out<=0;
   8327: out<=0;
   8328: out<=0;
   8329: out<=0;
   8330: out<=0;
   8331: out<=0;
   8332: out<=1;
   8333: out<=0;
   8334: out<=0;
   8335: out<=1;
   8336: out<=0;
   8337: out<=0;
   8338: out<=1;
   8339: out<=1;
   8340: out<=0;
   8341: out<=1;
   8342: out<=0;
   8343: out<=1;
   8344: out<=1;
   8345: out<=0;
   8346: out<=0;
   8347: out<=1;
   8348: out<=1;
   8349: out<=1;
   8350: out<=1;
   8351: out<=1;
   8352: out<=0;
   8353: out<=0;
   8354: out<=0;
   8355: out<=0;
   8356: out<=0;
   8357: out<=1;
   8358: out<=1;
   8359: out<=0;
   8360: out<=0;
   8361: out<=1;
   8362: out<=0;
   8363: out<=1;
   8364: out<=0;
   8365: out<=0;
   8366: out<=1;
   8367: out<=1;
   8368: out<=0;
   8369: out<=1;
   8370: out<=1;
   8371: out<=0;
   8372: out<=1;
   8373: out<=1;
   8374: out<=1;
   8375: out<=1;
   8376: out<=1;
   8377: out<=1;
   8378: out<=0;
   8379: out<=0;
   8380: out<=0;
   8381: out<=1;
   8382: out<=0;
   8383: out<=1;
   8384: out<=1;
   8385: out<=0;
   8386: out<=1;
   8387: out<=0;
   8388: out<=0;
   8389: out<=0;
   8390: out<=1;
   8391: out<=1;
   8392: out<=1;
   8393: out<=1;
   8394: out<=1;
   8395: out<=1;
   8396: out<=0;
   8397: out<=1;
   8398: out<=1;
   8399: out<=0;
   8400: out<=0;
   8401: out<=0;
   8402: out<=1;
   8403: out<=1;
   8404: out<=0;
   8405: out<=1;
   8406: out<=0;
   8407: out<=1;
   8408: out<=1;
   8409: out<=0;
   8410: out<=0;
   8411: out<=1;
   8412: out<=1;
   8413: out<=1;
   8414: out<=1;
   8415: out<=1;
   8416: out<=0;
   8417: out<=0;
   8418: out<=0;
   8419: out<=0;
   8420: out<=0;
   8421: out<=1;
   8422: out<=1;
   8423: out<=0;
   8424: out<=0;
   8425: out<=1;
   8426: out<=0;
   8427: out<=1;
   8428: out<=0;
   8429: out<=0;
   8430: out<=1;
   8431: out<=1;
   8432: out<=1;
   8433: out<=0;
   8434: out<=0;
   8435: out<=1;
   8436: out<=0;
   8437: out<=0;
   8438: out<=0;
   8439: out<=0;
   8440: out<=0;
   8441: out<=0;
   8442: out<=1;
   8443: out<=1;
   8444: out<=1;
   8445: out<=0;
   8446: out<=1;
   8447: out<=0;
   8448: out<=1;
   8449: out<=1;
   8450: out<=0;
   8451: out<=0;
   8452: out<=1;
   8453: out<=0;
   8454: out<=1;
   8455: out<=0;
   8456: out<=0;
   8457: out<=1;
   8458: out<=1;
   8459: out<=0;
   8460: out<=0;
   8461: out<=0;
   8462: out<=0;
   8463: out<=0;
   8464: out<=1;
   8465: out<=0;
   8466: out<=1;
   8467: out<=0;
   8468: out<=0;
   8469: out<=0;
   8470: out<=1;
   8471: out<=1;
   8472: out<=1;
   8473: out<=1;
   8474: out<=1;
   8475: out<=1;
   8476: out<=0;
   8477: out<=1;
   8478: out<=1;
   8479: out<=0;
   8480: out<=0;
   8481: out<=1;
   8482: out<=1;
   8483: out<=0;
   8484: out<=1;
   8485: out<=1;
   8486: out<=1;
   8487: out<=1;
   8488: out<=1;
   8489: out<=1;
   8490: out<=0;
   8491: out<=0;
   8492: out<=0;
   8493: out<=1;
   8494: out<=0;
   8495: out<=1;
   8496: out<=0;
   8497: out<=0;
   8498: out<=0;
   8499: out<=0;
   8500: out<=0;
   8501: out<=1;
   8502: out<=1;
   8503: out<=0;
   8504: out<=0;
   8505: out<=1;
   8506: out<=0;
   8507: out<=1;
   8508: out<=0;
   8509: out<=0;
   8510: out<=1;
   8511: out<=1;
   8512: out<=1;
   8513: out<=1;
   8514: out<=0;
   8515: out<=0;
   8516: out<=1;
   8517: out<=0;
   8518: out<=1;
   8519: out<=0;
   8520: out<=0;
   8521: out<=1;
   8522: out<=1;
   8523: out<=0;
   8524: out<=0;
   8525: out<=0;
   8526: out<=0;
   8527: out<=0;
   8528: out<=0;
   8529: out<=1;
   8530: out<=0;
   8531: out<=1;
   8532: out<=1;
   8533: out<=1;
   8534: out<=0;
   8535: out<=0;
   8536: out<=0;
   8537: out<=0;
   8538: out<=0;
   8539: out<=0;
   8540: out<=1;
   8541: out<=0;
   8542: out<=0;
   8543: out<=1;
   8544: out<=1;
   8545: out<=0;
   8546: out<=0;
   8547: out<=1;
   8548: out<=0;
   8549: out<=0;
   8550: out<=0;
   8551: out<=0;
   8552: out<=0;
   8553: out<=0;
   8554: out<=1;
   8555: out<=1;
   8556: out<=1;
   8557: out<=0;
   8558: out<=1;
   8559: out<=0;
   8560: out<=0;
   8561: out<=0;
   8562: out<=0;
   8563: out<=0;
   8564: out<=0;
   8565: out<=1;
   8566: out<=1;
   8567: out<=0;
   8568: out<=0;
   8569: out<=1;
   8570: out<=0;
   8571: out<=1;
   8572: out<=0;
   8573: out<=0;
   8574: out<=1;
   8575: out<=1;
   8576: out<=0;
   8577: out<=0;
   8578: out<=1;
   8579: out<=1;
   8580: out<=0;
   8581: out<=1;
   8582: out<=0;
   8583: out<=1;
   8584: out<=1;
   8585: out<=0;
   8586: out<=0;
   8587: out<=1;
   8588: out<=1;
   8589: out<=1;
   8590: out<=1;
   8591: out<=1;
   8592: out<=1;
   8593: out<=0;
   8594: out<=1;
   8595: out<=0;
   8596: out<=0;
   8597: out<=0;
   8598: out<=1;
   8599: out<=1;
   8600: out<=1;
   8601: out<=1;
   8602: out<=1;
   8603: out<=1;
   8604: out<=0;
   8605: out<=1;
   8606: out<=1;
   8607: out<=0;
   8608: out<=1;
   8609: out<=0;
   8610: out<=0;
   8611: out<=1;
   8612: out<=0;
   8613: out<=0;
   8614: out<=0;
   8615: out<=0;
   8616: out<=0;
   8617: out<=0;
   8618: out<=1;
   8619: out<=1;
   8620: out<=1;
   8621: out<=0;
   8622: out<=1;
   8623: out<=0;
   8624: out<=0;
   8625: out<=0;
   8626: out<=0;
   8627: out<=0;
   8628: out<=0;
   8629: out<=1;
   8630: out<=1;
   8631: out<=0;
   8632: out<=0;
   8633: out<=1;
   8634: out<=0;
   8635: out<=1;
   8636: out<=0;
   8637: out<=0;
   8638: out<=1;
   8639: out<=1;
   8640: out<=0;
   8641: out<=0;
   8642: out<=1;
   8643: out<=1;
   8644: out<=0;
   8645: out<=1;
   8646: out<=0;
   8647: out<=1;
   8648: out<=1;
   8649: out<=0;
   8650: out<=0;
   8651: out<=1;
   8652: out<=1;
   8653: out<=1;
   8654: out<=1;
   8655: out<=1;
   8656: out<=0;
   8657: out<=1;
   8658: out<=0;
   8659: out<=1;
   8660: out<=1;
   8661: out<=1;
   8662: out<=0;
   8663: out<=0;
   8664: out<=0;
   8665: out<=0;
   8666: out<=0;
   8667: out<=0;
   8668: out<=1;
   8669: out<=0;
   8670: out<=0;
   8671: out<=1;
   8672: out<=0;
   8673: out<=1;
   8674: out<=1;
   8675: out<=0;
   8676: out<=1;
   8677: out<=1;
   8678: out<=1;
   8679: out<=1;
   8680: out<=1;
   8681: out<=1;
   8682: out<=0;
   8683: out<=0;
   8684: out<=0;
   8685: out<=1;
   8686: out<=0;
   8687: out<=1;
   8688: out<=0;
   8689: out<=0;
   8690: out<=0;
   8691: out<=0;
   8692: out<=0;
   8693: out<=1;
   8694: out<=1;
   8695: out<=0;
   8696: out<=0;
   8697: out<=1;
   8698: out<=0;
   8699: out<=1;
   8700: out<=0;
   8701: out<=0;
   8702: out<=1;
   8703: out<=1;
   8704: out<=0;
   8705: out<=0;
   8706: out<=0;
   8707: out<=0;
   8708: out<=0;
   8709: out<=1;
   8710: out<=1;
   8711: out<=0;
   8712: out<=0;
   8713: out<=1;
   8714: out<=0;
   8715: out<=1;
   8716: out<=0;
   8717: out<=0;
   8718: out<=1;
   8719: out<=1;
   8720: out<=0;
   8721: out<=1;
   8722: out<=1;
   8723: out<=0;
   8724: out<=1;
   8725: out<=1;
   8726: out<=1;
   8727: out<=1;
   8728: out<=1;
   8729: out<=1;
   8730: out<=0;
   8731: out<=0;
   8732: out<=0;
   8733: out<=1;
   8734: out<=0;
   8735: out<=1;
   8736: out<=0;
   8737: out<=1;
   8738: out<=0;
   8739: out<=1;
   8740: out<=1;
   8741: out<=1;
   8742: out<=0;
   8743: out<=0;
   8744: out<=0;
   8745: out<=0;
   8746: out<=0;
   8747: out<=0;
   8748: out<=1;
   8749: out<=0;
   8750: out<=0;
   8751: out<=1;
   8752: out<=0;
   8753: out<=0;
   8754: out<=1;
   8755: out<=1;
   8756: out<=0;
   8757: out<=1;
   8758: out<=0;
   8759: out<=1;
   8760: out<=1;
   8761: out<=0;
   8762: out<=0;
   8763: out<=1;
   8764: out<=1;
   8765: out<=1;
   8766: out<=1;
   8767: out<=1;
   8768: out<=0;
   8769: out<=0;
   8770: out<=0;
   8771: out<=0;
   8772: out<=0;
   8773: out<=1;
   8774: out<=1;
   8775: out<=0;
   8776: out<=0;
   8777: out<=1;
   8778: out<=0;
   8779: out<=1;
   8780: out<=0;
   8781: out<=0;
   8782: out<=1;
   8783: out<=1;
   8784: out<=1;
   8785: out<=0;
   8786: out<=0;
   8787: out<=1;
   8788: out<=0;
   8789: out<=0;
   8790: out<=0;
   8791: out<=0;
   8792: out<=0;
   8793: out<=0;
   8794: out<=1;
   8795: out<=1;
   8796: out<=1;
   8797: out<=0;
   8798: out<=1;
   8799: out<=0;
   8800: out<=1;
   8801: out<=0;
   8802: out<=1;
   8803: out<=0;
   8804: out<=0;
   8805: out<=0;
   8806: out<=1;
   8807: out<=1;
   8808: out<=1;
   8809: out<=1;
   8810: out<=1;
   8811: out<=1;
   8812: out<=0;
   8813: out<=1;
   8814: out<=1;
   8815: out<=0;
   8816: out<=0;
   8817: out<=0;
   8818: out<=1;
   8819: out<=1;
   8820: out<=0;
   8821: out<=1;
   8822: out<=0;
   8823: out<=1;
   8824: out<=1;
   8825: out<=0;
   8826: out<=0;
   8827: out<=1;
   8828: out<=1;
   8829: out<=1;
   8830: out<=1;
   8831: out<=1;
   8832: out<=0;
   8833: out<=0;
   8834: out<=0;
   8835: out<=0;
   8836: out<=0;
   8837: out<=1;
   8838: out<=1;
   8839: out<=0;
   8840: out<=0;
   8841: out<=1;
   8842: out<=0;
   8843: out<=1;
   8844: out<=0;
   8845: out<=0;
   8846: out<=1;
   8847: out<=1;
   8848: out<=1;
   8849: out<=0;
   8850: out<=0;
   8851: out<=1;
   8852: out<=0;
   8853: out<=0;
   8854: out<=0;
   8855: out<=0;
   8856: out<=0;
   8857: out<=0;
   8858: out<=1;
   8859: out<=1;
   8860: out<=1;
   8861: out<=0;
   8862: out<=1;
   8863: out<=0;
   8864: out<=0;
   8865: out<=1;
   8866: out<=0;
   8867: out<=1;
   8868: out<=1;
   8869: out<=1;
   8870: out<=0;
   8871: out<=0;
   8872: out<=0;
   8873: out<=0;
   8874: out<=0;
   8875: out<=0;
   8876: out<=1;
   8877: out<=0;
   8878: out<=0;
   8879: out<=1;
   8880: out<=1;
   8881: out<=1;
   8882: out<=0;
   8883: out<=0;
   8884: out<=1;
   8885: out<=0;
   8886: out<=1;
   8887: out<=0;
   8888: out<=0;
   8889: out<=1;
   8890: out<=1;
   8891: out<=0;
   8892: out<=0;
   8893: out<=0;
   8894: out<=0;
   8895: out<=0;
   8896: out<=0;
   8897: out<=0;
   8898: out<=0;
   8899: out<=0;
   8900: out<=0;
   8901: out<=1;
   8902: out<=1;
   8903: out<=0;
   8904: out<=0;
   8905: out<=1;
   8906: out<=0;
   8907: out<=1;
   8908: out<=0;
   8909: out<=0;
   8910: out<=1;
   8911: out<=1;
   8912: out<=0;
   8913: out<=1;
   8914: out<=1;
   8915: out<=0;
   8916: out<=1;
   8917: out<=1;
   8918: out<=1;
   8919: out<=1;
   8920: out<=1;
   8921: out<=1;
   8922: out<=0;
   8923: out<=0;
   8924: out<=0;
   8925: out<=1;
   8926: out<=0;
   8927: out<=1;
   8928: out<=1;
   8929: out<=0;
   8930: out<=1;
   8931: out<=0;
   8932: out<=0;
   8933: out<=0;
   8934: out<=1;
   8935: out<=1;
   8936: out<=1;
   8937: out<=1;
   8938: out<=1;
   8939: out<=1;
   8940: out<=0;
   8941: out<=1;
   8942: out<=1;
   8943: out<=0;
   8944: out<=1;
   8945: out<=1;
   8946: out<=0;
   8947: out<=0;
   8948: out<=1;
   8949: out<=0;
   8950: out<=1;
   8951: out<=0;
   8952: out<=0;
   8953: out<=1;
   8954: out<=1;
   8955: out<=0;
   8956: out<=0;
   8957: out<=0;
   8958: out<=0;
   8959: out<=0;
   8960: out<=1;
   8961: out<=0;
   8962: out<=0;
   8963: out<=1;
   8964: out<=0;
   8965: out<=0;
   8966: out<=0;
   8967: out<=0;
   8968: out<=0;
   8969: out<=0;
   8970: out<=1;
   8971: out<=1;
   8972: out<=1;
   8973: out<=0;
   8974: out<=1;
   8975: out<=0;
   8976: out<=0;
   8977: out<=0;
   8978: out<=0;
   8979: out<=0;
   8980: out<=0;
   8981: out<=1;
   8982: out<=1;
   8983: out<=0;
   8984: out<=0;
   8985: out<=1;
   8986: out<=0;
   8987: out<=1;
   8988: out<=0;
   8989: out<=0;
   8990: out<=1;
   8991: out<=1;
   8992: out<=0;
   8993: out<=0;
   8994: out<=1;
   8995: out<=1;
   8996: out<=0;
   8997: out<=1;
   8998: out<=0;
   8999: out<=1;
   9000: out<=1;
   9001: out<=0;
   9002: out<=0;
   9003: out<=1;
   9004: out<=1;
   9005: out<=1;
   9006: out<=1;
   9007: out<=1;
   9008: out<=1;
   9009: out<=0;
   9010: out<=1;
   9011: out<=0;
   9012: out<=0;
   9013: out<=0;
   9014: out<=1;
   9015: out<=1;
   9016: out<=1;
   9017: out<=1;
   9018: out<=1;
   9019: out<=1;
   9020: out<=0;
   9021: out<=1;
   9022: out<=1;
   9023: out<=0;
   9024: out<=0;
   9025: out<=1;
   9026: out<=1;
   9027: out<=0;
   9028: out<=1;
   9029: out<=1;
   9030: out<=1;
   9031: out<=1;
   9032: out<=1;
   9033: out<=1;
   9034: out<=0;
   9035: out<=0;
   9036: out<=0;
   9037: out<=1;
   9038: out<=0;
   9039: out<=1;
   9040: out<=0;
   9041: out<=0;
   9042: out<=0;
   9043: out<=0;
   9044: out<=0;
   9045: out<=1;
   9046: out<=1;
   9047: out<=0;
   9048: out<=0;
   9049: out<=1;
   9050: out<=0;
   9051: out<=1;
   9052: out<=0;
   9053: out<=0;
   9054: out<=1;
   9055: out<=1;
   9056: out<=0;
   9057: out<=0;
   9058: out<=1;
   9059: out<=1;
   9060: out<=0;
   9061: out<=1;
   9062: out<=0;
   9063: out<=1;
   9064: out<=1;
   9065: out<=0;
   9066: out<=0;
   9067: out<=1;
   9068: out<=1;
   9069: out<=1;
   9070: out<=1;
   9071: out<=1;
   9072: out<=0;
   9073: out<=1;
   9074: out<=0;
   9075: out<=1;
   9076: out<=1;
   9077: out<=1;
   9078: out<=0;
   9079: out<=0;
   9080: out<=0;
   9081: out<=0;
   9082: out<=0;
   9083: out<=0;
   9084: out<=1;
   9085: out<=0;
   9086: out<=0;
   9087: out<=1;
   9088: out<=0;
   9089: out<=1;
   9090: out<=1;
   9091: out<=0;
   9092: out<=1;
   9093: out<=1;
   9094: out<=1;
   9095: out<=1;
   9096: out<=1;
   9097: out<=1;
   9098: out<=0;
   9099: out<=0;
   9100: out<=0;
   9101: out<=1;
   9102: out<=0;
   9103: out<=1;
   9104: out<=0;
   9105: out<=0;
   9106: out<=0;
   9107: out<=0;
   9108: out<=0;
   9109: out<=1;
   9110: out<=1;
   9111: out<=0;
   9112: out<=0;
   9113: out<=1;
   9114: out<=0;
   9115: out<=1;
   9116: out<=0;
   9117: out<=0;
   9118: out<=1;
   9119: out<=1;
   9120: out<=1;
   9121: out<=1;
   9122: out<=0;
   9123: out<=0;
   9124: out<=1;
   9125: out<=0;
   9126: out<=1;
   9127: out<=0;
   9128: out<=0;
   9129: out<=1;
   9130: out<=1;
   9131: out<=0;
   9132: out<=0;
   9133: out<=0;
   9134: out<=0;
   9135: out<=0;
   9136: out<=1;
   9137: out<=0;
   9138: out<=1;
   9139: out<=0;
   9140: out<=0;
   9141: out<=0;
   9142: out<=1;
   9143: out<=1;
   9144: out<=1;
   9145: out<=1;
   9146: out<=1;
   9147: out<=1;
   9148: out<=0;
   9149: out<=1;
   9150: out<=1;
   9151: out<=0;
   9152: out<=1;
   9153: out<=0;
   9154: out<=0;
   9155: out<=1;
   9156: out<=0;
   9157: out<=0;
   9158: out<=0;
   9159: out<=0;
   9160: out<=0;
   9161: out<=0;
   9162: out<=1;
   9163: out<=1;
   9164: out<=1;
   9165: out<=0;
   9166: out<=1;
   9167: out<=0;
   9168: out<=0;
   9169: out<=0;
   9170: out<=0;
   9171: out<=0;
   9172: out<=0;
   9173: out<=1;
   9174: out<=1;
   9175: out<=0;
   9176: out<=0;
   9177: out<=1;
   9178: out<=0;
   9179: out<=1;
   9180: out<=0;
   9181: out<=0;
   9182: out<=1;
   9183: out<=1;
   9184: out<=1;
   9185: out<=1;
   9186: out<=0;
   9187: out<=0;
   9188: out<=1;
   9189: out<=0;
   9190: out<=1;
   9191: out<=0;
   9192: out<=0;
   9193: out<=1;
   9194: out<=1;
   9195: out<=0;
   9196: out<=0;
   9197: out<=0;
   9198: out<=0;
   9199: out<=0;
   9200: out<=0;
   9201: out<=1;
   9202: out<=0;
   9203: out<=1;
   9204: out<=1;
   9205: out<=1;
   9206: out<=0;
   9207: out<=0;
   9208: out<=0;
   9209: out<=0;
   9210: out<=0;
   9211: out<=0;
   9212: out<=1;
   9213: out<=0;
   9214: out<=0;
   9215: out<=1;
   9216: out<=1;
   9217: out<=1;
   9218: out<=0;
   9219: out<=0;
   9220: out<=0;
   9221: out<=1;
   9222: out<=0;
   9223: out<=1;
   9224: out<=1;
   9225: out<=0;
   9226: out<=0;
   9227: out<=1;
   9228: out<=0;
   9229: out<=0;
   9230: out<=0;
   9231: out<=0;
   9232: out<=0;
   9233: out<=1;
   9234: out<=0;
   9235: out<=1;
   9236: out<=0;
   9237: out<=0;
   9238: out<=1;
   9239: out<=1;
   9240: out<=1;
   9241: out<=1;
   9242: out<=1;
   9243: out<=1;
   9244: out<=1;
   9245: out<=0;
   9246: out<=0;
   9247: out<=1;
   9248: out<=1;
   9249: out<=0;
   9250: out<=0;
   9251: out<=1;
   9252: out<=1;
   9253: out<=1;
   9254: out<=1;
   9255: out<=1;
   9256: out<=1;
   9257: out<=1;
   9258: out<=0;
   9259: out<=0;
   9260: out<=1;
   9261: out<=0;
   9262: out<=1;
   9263: out<=0;
   9264: out<=0;
   9265: out<=0;
   9266: out<=0;
   9267: out<=0;
   9268: out<=1;
   9269: out<=0;
   9270: out<=0;
   9271: out<=1;
   9272: out<=1;
   9273: out<=0;
   9274: out<=1;
   9275: out<=0;
   9276: out<=0;
   9277: out<=0;
   9278: out<=1;
   9279: out<=1;
   9280: out<=1;
   9281: out<=1;
   9282: out<=0;
   9283: out<=0;
   9284: out<=0;
   9285: out<=1;
   9286: out<=0;
   9287: out<=1;
   9288: out<=1;
   9289: out<=0;
   9290: out<=0;
   9291: out<=1;
   9292: out<=0;
   9293: out<=0;
   9294: out<=0;
   9295: out<=0;
   9296: out<=1;
   9297: out<=0;
   9298: out<=1;
   9299: out<=0;
   9300: out<=1;
   9301: out<=1;
   9302: out<=0;
   9303: out<=0;
   9304: out<=0;
   9305: out<=0;
   9306: out<=0;
   9307: out<=0;
   9308: out<=0;
   9309: out<=1;
   9310: out<=1;
   9311: out<=0;
   9312: out<=0;
   9313: out<=1;
   9314: out<=1;
   9315: out<=0;
   9316: out<=0;
   9317: out<=0;
   9318: out<=0;
   9319: out<=0;
   9320: out<=0;
   9321: out<=0;
   9322: out<=1;
   9323: out<=1;
   9324: out<=0;
   9325: out<=1;
   9326: out<=0;
   9327: out<=1;
   9328: out<=0;
   9329: out<=0;
   9330: out<=0;
   9331: out<=0;
   9332: out<=1;
   9333: out<=0;
   9334: out<=0;
   9335: out<=1;
   9336: out<=1;
   9337: out<=0;
   9338: out<=1;
   9339: out<=0;
   9340: out<=0;
   9341: out<=0;
   9342: out<=1;
   9343: out<=1;
   9344: out<=0;
   9345: out<=0;
   9346: out<=1;
   9347: out<=1;
   9348: out<=1;
   9349: out<=0;
   9350: out<=1;
   9351: out<=0;
   9352: out<=0;
   9353: out<=1;
   9354: out<=1;
   9355: out<=0;
   9356: out<=1;
   9357: out<=1;
   9358: out<=1;
   9359: out<=1;
   9360: out<=0;
   9361: out<=1;
   9362: out<=0;
   9363: out<=1;
   9364: out<=0;
   9365: out<=0;
   9366: out<=1;
   9367: out<=1;
   9368: out<=1;
   9369: out<=1;
   9370: out<=1;
   9371: out<=1;
   9372: out<=1;
   9373: out<=0;
   9374: out<=0;
   9375: out<=1;
   9376: out<=0;
   9377: out<=1;
   9378: out<=1;
   9379: out<=0;
   9380: out<=0;
   9381: out<=0;
   9382: out<=0;
   9383: out<=0;
   9384: out<=0;
   9385: out<=0;
   9386: out<=1;
   9387: out<=1;
   9388: out<=0;
   9389: out<=1;
   9390: out<=0;
   9391: out<=1;
   9392: out<=0;
   9393: out<=0;
   9394: out<=0;
   9395: out<=0;
   9396: out<=1;
   9397: out<=0;
   9398: out<=0;
   9399: out<=1;
   9400: out<=1;
   9401: out<=0;
   9402: out<=1;
   9403: out<=0;
   9404: out<=0;
   9405: out<=0;
   9406: out<=1;
   9407: out<=1;
   9408: out<=0;
   9409: out<=0;
   9410: out<=1;
   9411: out<=1;
   9412: out<=1;
   9413: out<=0;
   9414: out<=1;
   9415: out<=0;
   9416: out<=0;
   9417: out<=1;
   9418: out<=1;
   9419: out<=0;
   9420: out<=1;
   9421: out<=1;
   9422: out<=1;
   9423: out<=1;
   9424: out<=1;
   9425: out<=0;
   9426: out<=1;
   9427: out<=0;
   9428: out<=1;
   9429: out<=1;
   9430: out<=0;
   9431: out<=0;
   9432: out<=0;
   9433: out<=0;
   9434: out<=0;
   9435: out<=0;
   9436: out<=0;
   9437: out<=1;
   9438: out<=1;
   9439: out<=0;
   9440: out<=1;
   9441: out<=0;
   9442: out<=0;
   9443: out<=1;
   9444: out<=1;
   9445: out<=1;
   9446: out<=1;
   9447: out<=1;
   9448: out<=1;
   9449: out<=1;
   9450: out<=0;
   9451: out<=0;
   9452: out<=1;
   9453: out<=0;
   9454: out<=1;
   9455: out<=0;
   9456: out<=0;
   9457: out<=0;
   9458: out<=0;
   9459: out<=0;
   9460: out<=1;
   9461: out<=0;
   9462: out<=0;
   9463: out<=1;
   9464: out<=1;
   9465: out<=0;
   9466: out<=1;
   9467: out<=0;
   9468: out<=0;
   9469: out<=0;
   9470: out<=1;
   9471: out<=1;
   9472: out<=1;
   9473: out<=0;
   9474: out<=1;
   9475: out<=0;
   9476: out<=1;
   9477: out<=1;
   9478: out<=0;
   9479: out<=0;
   9480: out<=0;
   9481: out<=0;
   9482: out<=0;
   9483: out<=0;
   9484: out<=0;
   9485: out<=1;
   9486: out<=1;
   9487: out<=0;
   9488: out<=1;
   9489: out<=1;
   9490: out<=0;
   9491: out<=0;
   9492: out<=0;
   9493: out<=1;
   9494: out<=0;
   9495: out<=1;
   9496: out<=1;
   9497: out<=0;
   9498: out<=0;
   9499: out<=1;
   9500: out<=0;
   9501: out<=0;
   9502: out<=0;
   9503: out<=0;
   9504: out<=0;
   9505: out<=0;
   9506: out<=0;
   9507: out<=0;
   9508: out<=1;
   9509: out<=0;
   9510: out<=0;
   9511: out<=1;
   9512: out<=1;
   9513: out<=0;
   9514: out<=1;
   9515: out<=0;
   9516: out<=0;
   9517: out<=0;
   9518: out<=1;
   9519: out<=1;
   9520: out<=0;
   9521: out<=1;
   9522: out<=1;
   9523: out<=0;
   9524: out<=0;
   9525: out<=0;
   9526: out<=0;
   9527: out<=0;
   9528: out<=0;
   9529: out<=0;
   9530: out<=1;
   9531: out<=1;
   9532: out<=0;
   9533: out<=1;
   9534: out<=0;
   9535: out<=1;
   9536: out<=0;
   9537: out<=1;
   9538: out<=0;
   9539: out<=1;
   9540: out<=0;
   9541: out<=0;
   9542: out<=1;
   9543: out<=1;
   9544: out<=1;
   9545: out<=1;
   9546: out<=1;
   9547: out<=1;
   9548: out<=1;
   9549: out<=0;
   9550: out<=0;
   9551: out<=1;
   9552: out<=1;
   9553: out<=1;
   9554: out<=0;
   9555: out<=0;
   9556: out<=0;
   9557: out<=1;
   9558: out<=0;
   9559: out<=1;
   9560: out<=1;
   9561: out<=0;
   9562: out<=0;
   9563: out<=1;
   9564: out<=0;
   9565: out<=0;
   9566: out<=0;
   9567: out<=0;
   9568: out<=0;
   9569: out<=0;
   9570: out<=0;
   9571: out<=0;
   9572: out<=1;
   9573: out<=0;
   9574: out<=0;
   9575: out<=1;
   9576: out<=1;
   9577: out<=0;
   9578: out<=1;
   9579: out<=0;
   9580: out<=0;
   9581: out<=0;
   9582: out<=1;
   9583: out<=1;
   9584: out<=1;
   9585: out<=0;
   9586: out<=0;
   9587: out<=1;
   9588: out<=1;
   9589: out<=1;
   9590: out<=1;
   9591: out<=1;
   9592: out<=1;
   9593: out<=1;
   9594: out<=0;
   9595: out<=0;
   9596: out<=1;
   9597: out<=0;
   9598: out<=1;
   9599: out<=0;
   9600: out<=1;
   9601: out<=0;
   9602: out<=1;
   9603: out<=0;
   9604: out<=1;
   9605: out<=1;
   9606: out<=0;
   9607: out<=0;
   9608: out<=0;
   9609: out<=0;
   9610: out<=0;
   9611: out<=0;
   9612: out<=0;
   9613: out<=1;
   9614: out<=1;
   9615: out<=0;
   9616: out<=0;
   9617: out<=0;
   9618: out<=1;
   9619: out<=1;
   9620: out<=1;
   9621: out<=0;
   9622: out<=1;
   9623: out<=0;
   9624: out<=0;
   9625: out<=1;
   9626: out<=1;
   9627: out<=0;
   9628: out<=1;
   9629: out<=1;
   9630: out<=1;
   9631: out<=1;
   9632: out<=0;
   9633: out<=0;
   9634: out<=0;
   9635: out<=0;
   9636: out<=1;
   9637: out<=0;
   9638: out<=0;
   9639: out<=1;
   9640: out<=1;
   9641: out<=0;
   9642: out<=1;
   9643: out<=0;
   9644: out<=0;
   9645: out<=0;
   9646: out<=1;
   9647: out<=1;
   9648: out<=1;
   9649: out<=0;
   9650: out<=0;
   9651: out<=1;
   9652: out<=1;
   9653: out<=1;
   9654: out<=1;
   9655: out<=1;
   9656: out<=1;
   9657: out<=1;
   9658: out<=0;
   9659: out<=0;
   9660: out<=1;
   9661: out<=0;
   9662: out<=1;
   9663: out<=0;
   9664: out<=0;
   9665: out<=1;
   9666: out<=0;
   9667: out<=1;
   9668: out<=0;
   9669: out<=0;
   9670: out<=1;
   9671: out<=1;
   9672: out<=1;
   9673: out<=1;
   9674: out<=1;
   9675: out<=1;
   9676: out<=1;
   9677: out<=0;
   9678: out<=0;
   9679: out<=1;
   9680: out<=0;
   9681: out<=0;
   9682: out<=1;
   9683: out<=1;
   9684: out<=1;
   9685: out<=0;
   9686: out<=1;
   9687: out<=0;
   9688: out<=0;
   9689: out<=1;
   9690: out<=1;
   9691: out<=0;
   9692: out<=1;
   9693: out<=1;
   9694: out<=1;
   9695: out<=1;
   9696: out<=0;
   9697: out<=0;
   9698: out<=0;
   9699: out<=0;
   9700: out<=1;
   9701: out<=0;
   9702: out<=0;
   9703: out<=1;
   9704: out<=1;
   9705: out<=0;
   9706: out<=1;
   9707: out<=0;
   9708: out<=0;
   9709: out<=0;
   9710: out<=1;
   9711: out<=1;
   9712: out<=0;
   9713: out<=1;
   9714: out<=1;
   9715: out<=0;
   9716: out<=0;
   9717: out<=0;
   9718: out<=0;
   9719: out<=0;
   9720: out<=0;
   9721: out<=0;
   9722: out<=1;
   9723: out<=1;
   9724: out<=0;
   9725: out<=1;
   9726: out<=0;
   9727: out<=1;
   9728: out<=0;
   9729: out<=1;
   9730: out<=1;
   9731: out<=0;
   9732: out<=0;
   9733: out<=0;
   9734: out<=0;
   9735: out<=0;
   9736: out<=0;
   9737: out<=0;
   9738: out<=1;
   9739: out<=1;
   9740: out<=0;
   9741: out<=1;
   9742: out<=0;
   9743: out<=1;
   9744: out<=0;
   9745: out<=0;
   9746: out<=0;
   9747: out<=0;
   9748: out<=1;
   9749: out<=0;
   9750: out<=0;
   9751: out<=1;
   9752: out<=1;
   9753: out<=0;
   9754: out<=1;
   9755: out<=0;
   9756: out<=0;
   9757: out<=0;
   9758: out<=1;
   9759: out<=1;
   9760: out<=0;
   9761: out<=0;
   9762: out<=1;
   9763: out<=1;
   9764: out<=1;
   9765: out<=0;
   9766: out<=1;
   9767: out<=0;
   9768: out<=0;
   9769: out<=1;
   9770: out<=1;
   9771: out<=0;
   9772: out<=1;
   9773: out<=1;
   9774: out<=1;
   9775: out<=1;
   9776: out<=0;
   9777: out<=1;
   9778: out<=0;
   9779: out<=1;
   9780: out<=0;
   9781: out<=0;
   9782: out<=1;
   9783: out<=1;
   9784: out<=1;
   9785: out<=1;
   9786: out<=1;
   9787: out<=1;
   9788: out<=1;
   9789: out<=0;
   9790: out<=0;
   9791: out<=1;
   9792: out<=1;
   9793: out<=0;
   9794: out<=0;
   9795: out<=1;
   9796: out<=1;
   9797: out<=1;
   9798: out<=1;
   9799: out<=1;
   9800: out<=1;
   9801: out<=1;
   9802: out<=0;
   9803: out<=0;
   9804: out<=1;
   9805: out<=0;
   9806: out<=1;
   9807: out<=0;
   9808: out<=0;
   9809: out<=0;
   9810: out<=0;
   9811: out<=0;
   9812: out<=1;
   9813: out<=0;
   9814: out<=0;
   9815: out<=1;
   9816: out<=1;
   9817: out<=0;
   9818: out<=1;
   9819: out<=0;
   9820: out<=0;
   9821: out<=0;
   9822: out<=1;
   9823: out<=1;
   9824: out<=0;
   9825: out<=0;
   9826: out<=1;
   9827: out<=1;
   9828: out<=1;
   9829: out<=0;
   9830: out<=1;
   9831: out<=0;
   9832: out<=0;
   9833: out<=1;
   9834: out<=1;
   9835: out<=0;
   9836: out<=1;
   9837: out<=1;
   9838: out<=1;
   9839: out<=1;
   9840: out<=1;
   9841: out<=0;
   9842: out<=1;
   9843: out<=0;
   9844: out<=1;
   9845: out<=1;
   9846: out<=0;
   9847: out<=0;
   9848: out<=0;
   9849: out<=0;
   9850: out<=0;
   9851: out<=0;
   9852: out<=0;
   9853: out<=1;
   9854: out<=1;
   9855: out<=0;
   9856: out<=1;
   9857: out<=0;
   9858: out<=0;
   9859: out<=1;
   9860: out<=1;
   9861: out<=1;
   9862: out<=1;
   9863: out<=1;
   9864: out<=1;
   9865: out<=1;
   9866: out<=0;
   9867: out<=0;
   9868: out<=1;
   9869: out<=0;
   9870: out<=1;
   9871: out<=0;
   9872: out<=0;
   9873: out<=0;
   9874: out<=0;
   9875: out<=0;
   9876: out<=1;
   9877: out<=0;
   9878: out<=0;
   9879: out<=1;
   9880: out<=1;
   9881: out<=0;
   9882: out<=1;
   9883: out<=0;
   9884: out<=0;
   9885: out<=0;
   9886: out<=1;
   9887: out<=1;
   9888: out<=1;
   9889: out<=1;
   9890: out<=0;
   9891: out<=0;
   9892: out<=0;
   9893: out<=1;
   9894: out<=0;
   9895: out<=1;
   9896: out<=1;
   9897: out<=0;
   9898: out<=0;
   9899: out<=1;
   9900: out<=0;
   9901: out<=0;
   9902: out<=0;
   9903: out<=0;
   9904: out<=0;
   9905: out<=1;
   9906: out<=0;
   9907: out<=1;
   9908: out<=0;
   9909: out<=0;
   9910: out<=1;
   9911: out<=1;
   9912: out<=1;
   9913: out<=1;
   9914: out<=1;
   9915: out<=1;
   9916: out<=1;
   9917: out<=0;
   9918: out<=0;
   9919: out<=1;
   9920: out<=0;
   9921: out<=1;
   9922: out<=1;
   9923: out<=0;
   9924: out<=0;
   9925: out<=0;
   9926: out<=0;
   9927: out<=0;
   9928: out<=0;
   9929: out<=0;
   9930: out<=1;
   9931: out<=1;
   9932: out<=0;
   9933: out<=1;
   9934: out<=0;
   9935: out<=1;
   9936: out<=0;
   9937: out<=0;
   9938: out<=0;
   9939: out<=0;
   9940: out<=1;
   9941: out<=0;
   9942: out<=0;
   9943: out<=1;
   9944: out<=1;
   9945: out<=0;
   9946: out<=1;
   9947: out<=0;
   9948: out<=0;
   9949: out<=0;
   9950: out<=1;
   9951: out<=1;
   9952: out<=1;
   9953: out<=1;
   9954: out<=0;
   9955: out<=0;
   9956: out<=0;
   9957: out<=1;
   9958: out<=0;
   9959: out<=1;
   9960: out<=1;
   9961: out<=0;
   9962: out<=0;
   9963: out<=1;
   9964: out<=0;
   9965: out<=0;
   9966: out<=0;
   9967: out<=0;
   9968: out<=1;
   9969: out<=0;
   9970: out<=1;
   9971: out<=0;
   9972: out<=1;
   9973: out<=1;
   9974: out<=0;
   9975: out<=0;
   9976: out<=0;
   9977: out<=0;
   9978: out<=0;
   9979: out<=0;
   9980: out<=0;
   9981: out<=1;
   9982: out<=1;
   9983: out<=0;
   9984: out<=0;
   9985: out<=0;
   9986: out<=0;
   9987: out<=0;
   9988: out<=1;
   9989: out<=0;
   9990: out<=0;
   9991: out<=1;
   9992: out<=1;
   9993: out<=0;
   9994: out<=1;
   9995: out<=0;
   9996: out<=0;
   9997: out<=0;
   9998: out<=1;
   9999: out<=1;
   10000: out<=1;
   10001: out<=0;
   10002: out<=0;
   10003: out<=1;
   10004: out<=1;
   10005: out<=1;
   10006: out<=1;
   10007: out<=1;
   10008: out<=1;
   10009: out<=1;
   10010: out<=0;
   10011: out<=0;
   10012: out<=1;
   10013: out<=0;
   10014: out<=1;
   10015: out<=0;
   10016: out<=1;
   10017: out<=0;
   10018: out<=1;
   10019: out<=0;
   10020: out<=1;
   10021: out<=1;
   10022: out<=0;
   10023: out<=0;
   10024: out<=0;
   10025: out<=0;
   10026: out<=0;
   10027: out<=0;
   10028: out<=0;
   10029: out<=1;
   10030: out<=1;
   10031: out<=0;
   10032: out<=0;
   10033: out<=0;
   10034: out<=1;
   10035: out<=1;
   10036: out<=1;
   10037: out<=0;
   10038: out<=1;
   10039: out<=0;
   10040: out<=0;
   10041: out<=1;
   10042: out<=1;
   10043: out<=0;
   10044: out<=1;
   10045: out<=1;
   10046: out<=1;
   10047: out<=1;
   10048: out<=0;
   10049: out<=0;
   10050: out<=0;
   10051: out<=0;
   10052: out<=1;
   10053: out<=0;
   10054: out<=0;
   10055: out<=1;
   10056: out<=1;
   10057: out<=0;
   10058: out<=1;
   10059: out<=0;
   10060: out<=0;
   10061: out<=0;
   10062: out<=1;
   10063: out<=1;
   10064: out<=0;
   10065: out<=1;
   10066: out<=1;
   10067: out<=0;
   10068: out<=0;
   10069: out<=0;
   10070: out<=0;
   10071: out<=0;
   10072: out<=0;
   10073: out<=0;
   10074: out<=1;
   10075: out<=1;
   10076: out<=0;
   10077: out<=1;
   10078: out<=0;
   10079: out<=1;
   10080: out<=0;
   10081: out<=1;
   10082: out<=0;
   10083: out<=1;
   10084: out<=0;
   10085: out<=0;
   10086: out<=1;
   10087: out<=1;
   10088: out<=1;
   10089: out<=1;
   10090: out<=1;
   10091: out<=1;
   10092: out<=1;
   10093: out<=0;
   10094: out<=0;
   10095: out<=1;
   10096: out<=0;
   10097: out<=0;
   10098: out<=1;
   10099: out<=1;
   10100: out<=1;
   10101: out<=0;
   10102: out<=1;
   10103: out<=0;
   10104: out<=0;
   10105: out<=1;
   10106: out<=1;
   10107: out<=0;
   10108: out<=1;
   10109: out<=1;
   10110: out<=1;
   10111: out<=1;
   10112: out<=0;
   10113: out<=0;
   10114: out<=0;
   10115: out<=0;
   10116: out<=1;
   10117: out<=0;
   10118: out<=0;
   10119: out<=1;
   10120: out<=1;
   10121: out<=0;
   10122: out<=1;
   10123: out<=0;
   10124: out<=0;
   10125: out<=0;
   10126: out<=1;
   10127: out<=1;
   10128: out<=0;
   10129: out<=1;
   10130: out<=1;
   10131: out<=0;
   10132: out<=0;
   10133: out<=0;
   10134: out<=0;
   10135: out<=0;
   10136: out<=0;
   10137: out<=0;
   10138: out<=1;
   10139: out<=1;
   10140: out<=0;
   10141: out<=1;
   10142: out<=0;
   10143: out<=1;
   10144: out<=1;
   10145: out<=0;
   10146: out<=1;
   10147: out<=0;
   10148: out<=1;
   10149: out<=1;
   10150: out<=0;
   10151: out<=0;
   10152: out<=0;
   10153: out<=0;
   10154: out<=0;
   10155: out<=0;
   10156: out<=0;
   10157: out<=1;
   10158: out<=1;
   10159: out<=0;
   10160: out<=1;
   10161: out<=1;
   10162: out<=0;
   10163: out<=0;
   10164: out<=0;
   10165: out<=1;
   10166: out<=0;
   10167: out<=1;
   10168: out<=1;
   10169: out<=0;
   10170: out<=0;
   10171: out<=1;
   10172: out<=0;
   10173: out<=0;
   10174: out<=0;
   10175: out<=0;
   10176: out<=0;
   10177: out<=0;
   10178: out<=0;
   10179: out<=0;
   10180: out<=1;
   10181: out<=0;
   10182: out<=0;
   10183: out<=1;
   10184: out<=1;
   10185: out<=0;
   10186: out<=1;
   10187: out<=0;
   10188: out<=0;
   10189: out<=0;
   10190: out<=1;
   10191: out<=1;
   10192: out<=1;
   10193: out<=0;
   10194: out<=0;
   10195: out<=1;
   10196: out<=1;
   10197: out<=1;
   10198: out<=1;
   10199: out<=1;
   10200: out<=1;
   10201: out<=1;
   10202: out<=0;
   10203: out<=0;
   10204: out<=1;
   10205: out<=0;
   10206: out<=1;
   10207: out<=0;
   10208: out<=0;
   10209: out<=1;
   10210: out<=0;
   10211: out<=1;
   10212: out<=0;
   10213: out<=0;
   10214: out<=1;
   10215: out<=1;
   10216: out<=1;
   10217: out<=1;
   10218: out<=1;
   10219: out<=1;
   10220: out<=1;
   10221: out<=0;
   10222: out<=0;
   10223: out<=1;
   10224: out<=1;
   10225: out<=1;
   10226: out<=0;
   10227: out<=0;
   10228: out<=0;
   10229: out<=1;
   10230: out<=0;
   10231: out<=1;
   10232: out<=1;
   10233: out<=0;
   10234: out<=0;
   10235: out<=1;
   10236: out<=0;
   10237: out<=0;
   10238: out<=0;
   10239: out<=0;
   10240: out<=0;
   10241: out<=0;
   10242: out<=0;
   10243: out<=0;
   10244: out<=1;
   10245: out<=0;
   10246: out<=0;
   10247: out<=1;
   10248: out<=0;
   10249: out<=1;
   10250: out<=0;
   10251: out<=1;
   10252: out<=1;
   10253: out<=1;
   10254: out<=0;
   10255: out<=0;
   10256: out<=1;
   10257: out<=0;
   10258: out<=0;
   10259: out<=1;
   10260: out<=1;
   10261: out<=1;
   10262: out<=1;
   10263: out<=1;
   10264: out<=0;
   10265: out<=0;
   10266: out<=1;
   10267: out<=1;
   10268: out<=0;
   10269: out<=1;
   10270: out<=0;
   10271: out<=1;
   10272: out<=0;
   10273: out<=1;
   10274: out<=0;
   10275: out<=1;
   10276: out<=0;
   10277: out<=0;
   10278: out<=1;
   10279: out<=1;
   10280: out<=0;
   10281: out<=0;
   10282: out<=0;
   10283: out<=0;
   10284: out<=0;
   10285: out<=1;
   10286: out<=1;
   10287: out<=0;
   10288: out<=1;
   10289: out<=1;
   10290: out<=0;
   10291: out<=0;
   10292: out<=0;
   10293: out<=1;
   10294: out<=0;
   10295: out<=1;
   10296: out<=0;
   10297: out<=1;
   10298: out<=1;
   10299: out<=0;
   10300: out<=1;
   10301: out<=1;
   10302: out<=1;
   10303: out<=1;
   10304: out<=0;
   10305: out<=0;
   10306: out<=0;
   10307: out<=0;
   10308: out<=1;
   10309: out<=0;
   10310: out<=0;
   10311: out<=1;
   10312: out<=0;
   10313: out<=1;
   10314: out<=0;
   10315: out<=1;
   10316: out<=1;
   10317: out<=1;
   10318: out<=0;
   10319: out<=0;
   10320: out<=0;
   10321: out<=1;
   10322: out<=1;
   10323: out<=0;
   10324: out<=0;
   10325: out<=0;
   10326: out<=0;
   10327: out<=0;
   10328: out<=1;
   10329: out<=1;
   10330: out<=0;
   10331: out<=0;
   10332: out<=1;
   10333: out<=0;
   10334: out<=1;
   10335: out<=0;
   10336: out<=1;
   10337: out<=0;
   10338: out<=1;
   10339: out<=0;
   10340: out<=1;
   10341: out<=1;
   10342: out<=0;
   10343: out<=0;
   10344: out<=1;
   10345: out<=1;
   10346: out<=1;
   10347: out<=1;
   10348: out<=1;
   10349: out<=0;
   10350: out<=0;
   10351: out<=1;
   10352: out<=1;
   10353: out<=1;
   10354: out<=0;
   10355: out<=0;
   10356: out<=0;
   10357: out<=1;
   10358: out<=0;
   10359: out<=1;
   10360: out<=0;
   10361: out<=1;
   10362: out<=1;
   10363: out<=0;
   10364: out<=1;
   10365: out<=1;
   10366: out<=1;
   10367: out<=1;
   10368: out<=0;
   10369: out<=0;
   10370: out<=0;
   10371: out<=0;
   10372: out<=1;
   10373: out<=0;
   10374: out<=0;
   10375: out<=1;
   10376: out<=0;
   10377: out<=1;
   10378: out<=0;
   10379: out<=1;
   10380: out<=1;
   10381: out<=1;
   10382: out<=0;
   10383: out<=0;
   10384: out<=0;
   10385: out<=1;
   10386: out<=1;
   10387: out<=0;
   10388: out<=0;
   10389: out<=0;
   10390: out<=0;
   10391: out<=0;
   10392: out<=1;
   10393: out<=1;
   10394: out<=0;
   10395: out<=0;
   10396: out<=1;
   10397: out<=0;
   10398: out<=1;
   10399: out<=0;
   10400: out<=0;
   10401: out<=1;
   10402: out<=0;
   10403: out<=1;
   10404: out<=0;
   10405: out<=0;
   10406: out<=1;
   10407: out<=1;
   10408: out<=0;
   10409: out<=0;
   10410: out<=0;
   10411: out<=0;
   10412: out<=0;
   10413: out<=1;
   10414: out<=1;
   10415: out<=0;
   10416: out<=0;
   10417: out<=0;
   10418: out<=1;
   10419: out<=1;
   10420: out<=1;
   10421: out<=0;
   10422: out<=1;
   10423: out<=0;
   10424: out<=1;
   10425: out<=0;
   10426: out<=0;
   10427: out<=1;
   10428: out<=0;
   10429: out<=0;
   10430: out<=0;
   10431: out<=0;
   10432: out<=0;
   10433: out<=0;
   10434: out<=0;
   10435: out<=0;
   10436: out<=1;
   10437: out<=0;
   10438: out<=0;
   10439: out<=1;
   10440: out<=0;
   10441: out<=1;
   10442: out<=0;
   10443: out<=1;
   10444: out<=1;
   10445: out<=1;
   10446: out<=0;
   10447: out<=0;
   10448: out<=1;
   10449: out<=0;
   10450: out<=0;
   10451: out<=1;
   10452: out<=1;
   10453: out<=1;
   10454: out<=1;
   10455: out<=1;
   10456: out<=0;
   10457: out<=0;
   10458: out<=1;
   10459: out<=1;
   10460: out<=0;
   10461: out<=1;
   10462: out<=0;
   10463: out<=1;
   10464: out<=1;
   10465: out<=0;
   10466: out<=1;
   10467: out<=0;
   10468: out<=1;
   10469: out<=1;
   10470: out<=0;
   10471: out<=0;
   10472: out<=1;
   10473: out<=1;
   10474: out<=1;
   10475: out<=1;
   10476: out<=1;
   10477: out<=0;
   10478: out<=0;
   10479: out<=1;
   10480: out<=0;
   10481: out<=0;
   10482: out<=1;
   10483: out<=1;
   10484: out<=1;
   10485: out<=0;
   10486: out<=1;
   10487: out<=0;
   10488: out<=1;
   10489: out<=0;
   10490: out<=0;
   10491: out<=1;
   10492: out<=0;
   10493: out<=0;
   10494: out<=0;
   10495: out<=0;
   10496: out<=0;
   10497: out<=1;
   10498: out<=1;
   10499: out<=0;
   10500: out<=0;
   10501: out<=0;
   10502: out<=0;
   10503: out<=0;
   10504: out<=1;
   10505: out<=1;
   10506: out<=0;
   10507: out<=0;
   10508: out<=1;
   10509: out<=0;
   10510: out<=1;
   10511: out<=0;
   10512: out<=0;
   10513: out<=0;
   10514: out<=0;
   10515: out<=0;
   10516: out<=1;
   10517: out<=0;
   10518: out<=0;
   10519: out<=1;
   10520: out<=0;
   10521: out<=1;
   10522: out<=0;
   10523: out<=1;
   10524: out<=1;
   10525: out<=1;
   10526: out<=0;
   10527: out<=0;
   10528: out<=1;
   10529: out<=1;
   10530: out<=0;
   10531: out<=0;
   10532: out<=0;
   10533: out<=1;
   10534: out<=0;
   10535: out<=1;
   10536: out<=0;
   10537: out<=1;
   10538: out<=1;
   10539: out<=0;
   10540: out<=1;
   10541: out<=1;
   10542: out<=1;
   10543: out<=1;
   10544: out<=1;
   10545: out<=0;
   10546: out<=1;
   10547: out<=0;
   10548: out<=1;
   10549: out<=1;
   10550: out<=0;
   10551: out<=0;
   10552: out<=1;
   10553: out<=1;
   10554: out<=1;
   10555: out<=1;
   10556: out<=1;
   10557: out<=0;
   10558: out<=0;
   10559: out<=1;
   10560: out<=1;
   10561: out<=0;
   10562: out<=0;
   10563: out<=1;
   10564: out<=1;
   10565: out<=1;
   10566: out<=1;
   10567: out<=1;
   10568: out<=0;
   10569: out<=0;
   10570: out<=1;
   10571: out<=1;
   10572: out<=0;
   10573: out<=1;
   10574: out<=0;
   10575: out<=1;
   10576: out<=0;
   10577: out<=0;
   10578: out<=0;
   10579: out<=0;
   10580: out<=1;
   10581: out<=0;
   10582: out<=0;
   10583: out<=1;
   10584: out<=0;
   10585: out<=1;
   10586: out<=0;
   10587: out<=1;
   10588: out<=1;
   10589: out<=1;
   10590: out<=0;
   10591: out<=0;
   10592: out<=1;
   10593: out<=1;
   10594: out<=0;
   10595: out<=0;
   10596: out<=0;
   10597: out<=1;
   10598: out<=0;
   10599: out<=1;
   10600: out<=0;
   10601: out<=1;
   10602: out<=1;
   10603: out<=0;
   10604: out<=1;
   10605: out<=1;
   10606: out<=1;
   10607: out<=1;
   10608: out<=0;
   10609: out<=1;
   10610: out<=0;
   10611: out<=1;
   10612: out<=0;
   10613: out<=0;
   10614: out<=1;
   10615: out<=1;
   10616: out<=0;
   10617: out<=0;
   10618: out<=0;
   10619: out<=0;
   10620: out<=0;
   10621: out<=1;
   10622: out<=1;
   10623: out<=0;
   10624: out<=1;
   10625: out<=0;
   10626: out<=0;
   10627: out<=1;
   10628: out<=1;
   10629: out<=1;
   10630: out<=1;
   10631: out<=1;
   10632: out<=0;
   10633: out<=0;
   10634: out<=1;
   10635: out<=1;
   10636: out<=0;
   10637: out<=1;
   10638: out<=0;
   10639: out<=1;
   10640: out<=0;
   10641: out<=0;
   10642: out<=0;
   10643: out<=0;
   10644: out<=1;
   10645: out<=0;
   10646: out<=0;
   10647: out<=1;
   10648: out<=0;
   10649: out<=1;
   10650: out<=0;
   10651: out<=1;
   10652: out<=1;
   10653: out<=1;
   10654: out<=0;
   10655: out<=0;
   10656: out<=0;
   10657: out<=0;
   10658: out<=1;
   10659: out<=1;
   10660: out<=1;
   10661: out<=0;
   10662: out<=1;
   10663: out<=0;
   10664: out<=1;
   10665: out<=0;
   10666: out<=0;
   10667: out<=1;
   10668: out<=0;
   10669: out<=0;
   10670: out<=0;
   10671: out<=0;
   10672: out<=1;
   10673: out<=0;
   10674: out<=1;
   10675: out<=0;
   10676: out<=1;
   10677: out<=1;
   10678: out<=0;
   10679: out<=0;
   10680: out<=1;
   10681: out<=1;
   10682: out<=1;
   10683: out<=1;
   10684: out<=1;
   10685: out<=0;
   10686: out<=0;
   10687: out<=1;
   10688: out<=0;
   10689: out<=1;
   10690: out<=1;
   10691: out<=0;
   10692: out<=0;
   10693: out<=0;
   10694: out<=0;
   10695: out<=0;
   10696: out<=1;
   10697: out<=1;
   10698: out<=0;
   10699: out<=0;
   10700: out<=1;
   10701: out<=0;
   10702: out<=1;
   10703: out<=0;
   10704: out<=0;
   10705: out<=0;
   10706: out<=0;
   10707: out<=0;
   10708: out<=1;
   10709: out<=0;
   10710: out<=0;
   10711: out<=1;
   10712: out<=0;
   10713: out<=1;
   10714: out<=0;
   10715: out<=1;
   10716: out<=1;
   10717: out<=1;
   10718: out<=0;
   10719: out<=0;
   10720: out<=0;
   10721: out<=0;
   10722: out<=1;
   10723: out<=1;
   10724: out<=1;
   10725: out<=0;
   10726: out<=1;
   10727: out<=0;
   10728: out<=1;
   10729: out<=0;
   10730: out<=0;
   10731: out<=1;
   10732: out<=0;
   10733: out<=0;
   10734: out<=0;
   10735: out<=0;
   10736: out<=0;
   10737: out<=1;
   10738: out<=0;
   10739: out<=1;
   10740: out<=0;
   10741: out<=0;
   10742: out<=1;
   10743: out<=1;
   10744: out<=0;
   10745: out<=0;
   10746: out<=0;
   10747: out<=0;
   10748: out<=0;
   10749: out<=1;
   10750: out<=1;
   10751: out<=0;
   10752: out<=0;
   10753: out<=1;
   10754: out<=0;
   10755: out<=1;
   10756: out<=0;
   10757: out<=0;
   10758: out<=1;
   10759: out<=1;
   10760: out<=0;
   10761: out<=0;
   10762: out<=0;
   10763: out<=0;
   10764: out<=0;
   10765: out<=1;
   10766: out<=1;
   10767: out<=0;
   10768: out<=0;
   10769: out<=0;
   10770: out<=1;
   10771: out<=1;
   10772: out<=1;
   10773: out<=0;
   10774: out<=1;
   10775: out<=0;
   10776: out<=1;
   10777: out<=0;
   10778: out<=0;
   10779: out<=1;
   10780: out<=0;
   10781: out<=0;
   10782: out<=0;
   10783: out<=0;
   10784: out<=0;
   10785: out<=0;
   10786: out<=0;
   10787: out<=0;
   10788: out<=1;
   10789: out<=0;
   10790: out<=0;
   10791: out<=1;
   10792: out<=0;
   10793: out<=1;
   10794: out<=0;
   10795: out<=1;
   10796: out<=1;
   10797: out<=1;
   10798: out<=0;
   10799: out<=0;
   10800: out<=0;
   10801: out<=1;
   10802: out<=1;
   10803: out<=0;
   10804: out<=0;
   10805: out<=0;
   10806: out<=0;
   10807: out<=0;
   10808: out<=1;
   10809: out<=1;
   10810: out<=0;
   10811: out<=0;
   10812: out<=1;
   10813: out<=0;
   10814: out<=1;
   10815: out<=0;
   10816: out<=1;
   10817: out<=0;
   10818: out<=1;
   10819: out<=0;
   10820: out<=1;
   10821: out<=1;
   10822: out<=0;
   10823: out<=0;
   10824: out<=1;
   10825: out<=1;
   10826: out<=1;
   10827: out<=1;
   10828: out<=1;
   10829: out<=0;
   10830: out<=0;
   10831: out<=1;
   10832: out<=0;
   10833: out<=0;
   10834: out<=1;
   10835: out<=1;
   10836: out<=1;
   10837: out<=0;
   10838: out<=1;
   10839: out<=0;
   10840: out<=1;
   10841: out<=0;
   10842: out<=0;
   10843: out<=1;
   10844: out<=0;
   10845: out<=0;
   10846: out<=0;
   10847: out<=0;
   10848: out<=0;
   10849: out<=0;
   10850: out<=0;
   10851: out<=0;
   10852: out<=1;
   10853: out<=0;
   10854: out<=0;
   10855: out<=1;
   10856: out<=0;
   10857: out<=1;
   10858: out<=0;
   10859: out<=1;
   10860: out<=1;
   10861: out<=1;
   10862: out<=0;
   10863: out<=0;
   10864: out<=1;
   10865: out<=0;
   10866: out<=0;
   10867: out<=1;
   10868: out<=1;
   10869: out<=1;
   10870: out<=1;
   10871: out<=1;
   10872: out<=0;
   10873: out<=0;
   10874: out<=1;
   10875: out<=1;
   10876: out<=0;
   10877: out<=1;
   10878: out<=0;
   10879: out<=1;
   10880: out<=0;
   10881: out<=1;
   10882: out<=0;
   10883: out<=1;
   10884: out<=0;
   10885: out<=0;
   10886: out<=1;
   10887: out<=1;
   10888: out<=0;
   10889: out<=0;
   10890: out<=0;
   10891: out<=0;
   10892: out<=0;
   10893: out<=1;
   10894: out<=1;
   10895: out<=0;
   10896: out<=1;
   10897: out<=1;
   10898: out<=0;
   10899: out<=0;
   10900: out<=0;
   10901: out<=1;
   10902: out<=0;
   10903: out<=1;
   10904: out<=0;
   10905: out<=1;
   10906: out<=1;
   10907: out<=0;
   10908: out<=1;
   10909: out<=1;
   10910: out<=1;
   10911: out<=1;
   10912: out<=0;
   10913: out<=0;
   10914: out<=0;
   10915: out<=0;
   10916: out<=1;
   10917: out<=0;
   10918: out<=0;
   10919: out<=1;
   10920: out<=0;
   10921: out<=1;
   10922: out<=0;
   10923: out<=1;
   10924: out<=1;
   10925: out<=1;
   10926: out<=0;
   10927: out<=0;
   10928: out<=1;
   10929: out<=0;
   10930: out<=0;
   10931: out<=1;
   10932: out<=1;
   10933: out<=1;
   10934: out<=1;
   10935: out<=1;
   10936: out<=0;
   10937: out<=0;
   10938: out<=1;
   10939: out<=1;
   10940: out<=0;
   10941: out<=1;
   10942: out<=0;
   10943: out<=1;
   10944: out<=1;
   10945: out<=0;
   10946: out<=1;
   10947: out<=0;
   10948: out<=1;
   10949: out<=1;
   10950: out<=0;
   10951: out<=0;
   10952: out<=1;
   10953: out<=1;
   10954: out<=1;
   10955: out<=1;
   10956: out<=1;
   10957: out<=0;
   10958: out<=0;
   10959: out<=1;
   10960: out<=1;
   10961: out<=1;
   10962: out<=0;
   10963: out<=0;
   10964: out<=0;
   10965: out<=1;
   10966: out<=0;
   10967: out<=1;
   10968: out<=0;
   10969: out<=1;
   10970: out<=1;
   10971: out<=0;
   10972: out<=1;
   10973: out<=1;
   10974: out<=1;
   10975: out<=1;
   10976: out<=0;
   10977: out<=0;
   10978: out<=0;
   10979: out<=0;
   10980: out<=1;
   10981: out<=0;
   10982: out<=0;
   10983: out<=1;
   10984: out<=0;
   10985: out<=1;
   10986: out<=0;
   10987: out<=1;
   10988: out<=1;
   10989: out<=1;
   10990: out<=0;
   10991: out<=0;
   10992: out<=0;
   10993: out<=1;
   10994: out<=1;
   10995: out<=0;
   10996: out<=0;
   10997: out<=0;
   10998: out<=0;
   10999: out<=0;
   11000: out<=1;
   11001: out<=1;
   11002: out<=0;
   11003: out<=0;
   11004: out<=1;
   11005: out<=0;
   11006: out<=1;
   11007: out<=0;
   11008: out<=0;
   11009: out<=0;
   11010: out<=1;
   11011: out<=1;
   11012: out<=1;
   11013: out<=0;
   11014: out<=1;
   11015: out<=0;
   11016: out<=1;
   11017: out<=0;
   11018: out<=0;
   11019: out<=1;
   11020: out<=0;
   11021: out<=0;
   11022: out<=0;
   11023: out<=0;
   11024: out<=1;
   11025: out<=0;
   11026: out<=1;
   11027: out<=0;
   11028: out<=1;
   11029: out<=1;
   11030: out<=0;
   11031: out<=0;
   11032: out<=1;
   11033: out<=1;
   11034: out<=1;
   11035: out<=1;
   11036: out<=1;
   11037: out<=0;
   11038: out<=0;
   11039: out<=1;
   11040: out<=1;
   11041: out<=0;
   11042: out<=0;
   11043: out<=1;
   11044: out<=1;
   11045: out<=1;
   11046: out<=1;
   11047: out<=1;
   11048: out<=0;
   11049: out<=0;
   11050: out<=1;
   11051: out<=1;
   11052: out<=0;
   11053: out<=1;
   11054: out<=0;
   11055: out<=1;
   11056: out<=0;
   11057: out<=0;
   11058: out<=0;
   11059: out<=0;
   11060: out<=1;
   11061: out<=0;
   11062: out<=0;
   11063: out<=1;
   11064: out<=0;
   11065: out<=1;
   11066: out<=0;
   11067: out<=1;
   11068: out<=1;
   11069: out<=1;
   11070: out<=0;
   11071: out<=0;
   11072: out<=0;
   11073: out<=0;
   11074: out<=1;
   11075: out<=1;
   11076: out<=1;
   11077: out<=0;
   11078: out<=1;
   11079: out<=0;
   11080: out<=1;
   11081: out<=0;
   11082: out<=0;
   11083: out<=1;
   11084: out<=0;
   11085: out<=0;
   11086: out<=0;
   11087: out<=0;
   11088: out<=0;
   11089: out<=1;
   11090: out<=0;
   11091: out<=1;
   11092: out<=0;
   11093: out<=0;
   11094: out<=1;
   11095: out<=1;
   11096: out<=0;
   11097: out<=0;
   11098: out<=0;
   11099: out<=0;
   11100: out<=0;
   11101: out<=1;
   11102: out<=1;
   11103: out<=0;
   11104: out<=0;
   11105: out<=1;
   11106: out<=1;
   11107: out<=0;
   11108: out<=0;
   11109: out<=0;
   11110: out<=0;
   11111: out<=0;
   11112: out<=1;
   11113: out<=1;
   11114: out<=0;
   11115: out<=0;
   11116: out<=1;
   11117: out<=0;
   11118: out<=1;
   11119: out<=0;
   11120: out<=0;
   11121: out<=0;
   11122: out<=0;
   11123: out<=0;
   11124: out<=1;
   11125: out<=0;
   11126: out<=0;
   11127: out<=1;
   11128: out<=0;
   11129: out<=1;
   11130: out<=0;
   11131: out<=1;
   11132: out<=1;
   11133: out<=1;
   11134: out<=0;
   11135: out<=0;
   11136: out<=1;
   11137: out<=1;
   11138: out<=0;
   11139: out<=0;
   11140: out<=0;
   11141: out<=1;
   11142: out<=0;
   11143: out<=1;
   11144: out<=0;
   11145: out<=1;
   11146: out<=1;
   11147: out<=0;
   11148: out<=1;
   11149: out<=1;
   11150: out<=1;
   11151: out<=1;
   11152: out<=1;
   11153: out<=0;
   11154: out<=1;
   11155: out<=0;
   11156: out<=1;
   11157: out<=1;
   11158: out<=0;
   11159: out<=0;
   11160: out<=1;
   11161: out<=1;
   11162: out<=1;
   11163: out<=1;
   11164: out<=1;
   11165: out<=0;
   11166: out<=0;
   11167: out<=1;
   11168: out<=0;
   11169: out<=1;
   11170: out<=1;
   11171: out<=0;
   11172: out<=0;
   11173: out<=0;
   11174: out<=0;
   11175: out<=0;
   11176: out<=1;
   11177: out<=1;
   11178: out<=0;
   11179: out<=0;
   11180: out<=1;
   11181: out<=0;
   11182: out<=1;
   11183: out<=0;
   11184: out<=0;
   11185: out<=0;
   11186: out<=0;
   11187: out<=0;
   11188: out<=1;
   11189: out<=0;
   11190: out<=0;
   11191: out<=1;
   11192: out<=0;
   11193: out<=1;
   11194: out<=0;
   11195: out<=1;
   11196: out<=1;
   11197: out<=1;
   11198: out<=0;
   11199: out<=0;
   11200: out<=1;
   11201: out<=1;
   11202: out<=0;
   11203: out<=0;
   11204: out<=0;
   11205: out<=1;
   11206: out<=0;
   11207: out<=1;
   11208: out<=0;
   11209: out<=1;
   11210: out<=1;
   11211: out<=0;
   11212: out<=1;
   11213: out<=1;
   11214: out<=1;
   11215: out<=1;
   11216: out<=0;
   11217: out<=1;
   11218: out<=0;
   11219: out<=1;
   11220: out<=0;
   11221: out<=0;
   11222: out<=1;
   11223: out<=1;
   11224: out<=0;
   11225: out<=0;
   11226: out<=0;
   11227: out<=0;
   11228: out<=0;
   11229: out<=1;
   11230: out<=1;
   11231: out<=0;
   11232: out<=1;
   11233: out<=0;
   11234: out<=0;
   11235: out<=1;
   11236: out<=1;
   11237: out<=1;
   11238: out<=1;
   11239: out<=1;
   11240: out<=0;
   11241: out<=0;
   11242: out<=1;
   11243: out<=1;
   11244: out<=0;
   11245: out<=1;
   11246: out<=0;
   11247: out<=1;
   11248: out<=0;
   11249: out<=0;
   11250: out<=0;
   11251: out<=0;
   11252: out<=1;
   11253: out<=0;
   11254: out<=0;
   11255: out<=1;
   11256: out<=0;
   11257: out<=1;
   11258: out<=0;
   11259: out<=1;
   11260: out<=1;
   11261: out<=1;
   11262: out<=0;
   11263: out<=0;
   11264: out<=1;
   11265: out<=0;
   11266: out<=0;
   11267: out<=1;
   11268: out<=0;
   11269: out<=0;
   11270: out<=0;
   11271: out<=0;
   11272: out<=1;
   11273: out<=1;
   11274: out<=0;
   11275: out<=0;
   11276: out<=0;
   11277: out<=1;
   11278: out<=0;
   11279: out<=1;
   11280: out<=0;
   11281: out<=0;
   11282: out<=0;
   11283: out<=0;
   11284: out<=0;
   11285: out<=1;
   11286: out<=1;
   11287: out<=0;
   11288: out<=1;
   11289: out<=0;
   11290: out<=1;
   11291: out<=0;
   11292: out<=1;
   11293: out<=1;
   11294: out<=0;
   11295: out<=0;
   11296: out<=1;
   11297: out<=1;
   11298: out<=0;
   11299: out<=0;
   11300: out<=1;
   11301: out<=0;
   11302: out<=1;
   11303: out<=0;
   11304: out<=1;
   11305: out<=0;
   11306: out<=0;
   11307: out<=1;
   11308: out<=1;
   11309: out<=1;
   11310: out<=1;
   11311: out<=1;
   11312: out<=0;
   11313: out<=1;
   11314: out<=0;
   11315: out<=1;
   11316: out<=1;
   11317: out<=1;
   11318: out<=0;
   11319: out<=0;
   11320: out<=1;
   11321: out<=1;
   11322: out<=1;
   11323: out<=1;
   11324: out<=0;
   11325: out<=1;
   11326: out<=1;
   11327: out<=0;
   11328: out<=0;
   11329: out<=1;
   11330: out<=1;
   11331: out<=0;
   11332: out<=1;
   11333: out<=1;
   11334: out<=1;
   11335: out<=1;
   11336: out<=0;
   11337: out<=0;
   11338: out<=1;
   11339: out<=1;
   11340: out<=1;
   11341: out<=0;
   11342: out<=1;
   11343: out<=0;
   11344: out<=0;
   11345: out<=0;
   11346: out<=0;
   11347: out<=0;
   11348: out<=0;
   11349: out<=1;
   11350: out<=1;
   11351: out<=0;
   11352: out<=1;
   11353: out<=0;
   11354: out<=1;
   11355: out<=0;
   11356: out<=1;
   11357: out<=1;
   11358: out<=0;
   11359: out<=0;
   11360: out<=1;
   11361: out<=1;
   11362: out<=0;
   11363: out<=0;
   11364: out<=1;
   11365: out<=0;
   11366: out<=1;
   11367: out<=0;
   11368: out<=1;
   11369: out<=0;
   11370: out<=0;
   11371: out<=1;
   11372: out<=1;
   11373: out<=1;
   11374: out<=1;
   11375: out<=1;
   11376: out<=1;
   11377: out<=0;
   11378: out<=1;
   11379: out<=0;
   11380: out<=0;
   11381: out<=0;
   11382: out<=1;
   11383: out<=1;
   11384: out<=0;
   11385: out<=0;
   11386: out<=0;
   11387: out<=0;
   11388: out<=1;
   11389: out<=0;
   11390: out<=0;
   11391: out<=1;
   11392: out<=0;
   11393: out<=1;
   11394: out<=1;
   11395: out<=0;
   11396: out<=1;
   11397: out<=1;
   11398: out<=1;
   11399: out<=1;
   11400: out<=0;
   11401: out<=0;
   11402: out<=1;
   11403: out<=1;
   11404: out<=1;
   11405: out<=0;
   11406: out<=1;
   11407: out<=0;
   11408: out<=0;
   11409: out<=0;
   11410: out<=0;
   11411: out<=0;
   11412: out<=0;
   11413: out<=1;
   11414: out<=1;
   11415: out<=0;
   11416: out<=1;
   11417: out<=0;
   11418: out<=1;
   11419: out<=0;
   11420: out<=1;
   11421: out<=1;
   11422: out<=0;
   11423: out<=0;
   11424: out<=0;
   11425: out<=0;
   11426: out<=1;
   11427: out<=1;
   11428: out<=0;
   11429: out<=1;
   11430: out<=0;
   11431: out<=1;
   11432: out<=0;
   11433: out<=1;
   11434: out<=1;
   11435: out<=0;
   11436: out<=0;
   11437: out<=0;
   11438: out<=0;
   11439: out<=0;
   11440: out<=0;
   11441: out<=1;
   11442: out<=0;
   11443: out<=1;
   11444: out<=1;
   11445: out<=1;
   11446: out<=0;
   11447: out<=0;
   11448: out<=1;
   11449: out<=1;
   11450: out<=1;
   11451: out<=1;
   11452: out<=0;
   11453: out<=1;
   11454: out<=1;
   11455: out<=0;
   11456: out<=1;
   11457: out<=0;
   11458: out<=0;
   11459: out<=1;
   11460: out<=0;
   11461: out<=0;
   11462: out<=0;
   11463: out<=0;
   11464: out<=1;
   11465: out<=1;
   11466: out<=0;
   11467: out<=0;
   11468: out<=0;
   11469: out<=1;
   11470: out<=0;
   11471: out<=1;
   11472: out<=0;
   11473: out<=0;
   11474: out<=0;
   11475: out<=0;
   11476: out<=0;
   11477: out<=1;
   11478: out<=1;
   11479: out<=0;
   11480: out<=1;
   11481: out<=0;
   11482: out<=1;
   11483: out<=0;
   11484: out<=1;
   11485: out<=1;
   11486: out<=0;
   11487: out<=0;
   11488: out<=0;
   11489: out<=0;
   11490: out<=1;
   11491: out<=1;
   11492: out<=0;
   11493: out<=1;
   11494: out<=0;
   11495: out<=1;
   11496: out<=0;
   11497: out<=1;
   11498: out<=1;
   11499: out<=0;
   11500: out<=0;
   11501: out<=0;
   11502: out<=0;
   11503: out<=0;
   11504: out<=1;
   11505: out<=0;
   11506: out<=1;
   11507: out<=0;
   11508: out<=0;
   11509: out<=0;
   11510: out<=1;
   11511: out<=1;
   11512: out<=0;
   11513: out<=0;
   11514: out<=0;
   11515: out<=0;
   11516: out<=1;
   11517: out<=0;
   11518: out<=0;
   11519: out<=1;
   11520: out<=0;
   11521: out<=0;
   11522: out<=0;
   11523: out<=0;
   11524: out<=0;
   11525: out<=1;
   11526: out<=1;
   11527: out<=0;
   11528: out<=1;
   11529: out<=0;
   11530: out<=1;
   11531: out<=0;
   11532: out<=1;
   11533: out<=1;
   11534: out<=0;
   11535: out<=0;
   11536: out<=0;
   11537: out<=1;
   11538: out<=1;
   11539: out<=0;
   11540: out<=1;
   11541: out<=1;
   11542: out<=1;
   11543: out<=1;
   11544: out<=0;
   11545: out<=0;
   11546: out<=1;
   11547: out<=1;
   11548: out<=1;
   11549: out<=0;
   11550: out<=1;
   11551: out<=0;
   11552: out<=1;
   11553: out<=0;
   11554: out<=1;
   11555: out<=0;
   11556: out<=0;
   11557: out<=0;
   11558: out<=1;
   11559: out<=1;
   11560: out<=0;
   11561: out<=0;
   11562: out<=0;
   11563: out<=0;
   11564: out<=1;
   11565: out<=0;
   11566: out<=0;
   11567: out<=1;
   11568: out<=1;
   11569: out<=1;
   11570: out<=0;
   11571: out<=0;
   11572: out<=1;
   11573: out<=0;
   11574: out<=1;
   11575: out<=0;
   11576: out<=1;
   11577: out<=0;
   11578: out<=0;
   11579: out<=1;
   11580: out<=1;
   11581: out<=1;
   11582: out<=1;
   11583: out<=1;
   11584: out<=0;
   11585: out<=0;
   11586: out<=0;
   11587: out<=0;
   11588: out<=0;
   11589: out<=1;
   11590: out<=1;
   11591: out<=0;
   11592: out<=1;
   11593: out<=0;
   11594: out<=1;
   11595: out<=0;
   11596: out<=1;
   11597: out<=1;
   11598: out<=0;
   11599: out<=0;
   11600: out<=1;
   11601: out<=0;
   11602: out<=0;
   11603: out<=1;
   11604: out<=0;
   11605: out<=0;
   11606: out<=0;
   11607: out<=0;
   11608: out<=1;
   11609: out<=1;
   11610: out<=0;
   11611: out<=0;
   11612: out<=0;
   11613: out<=1;
   11614: out<=0;
   11615: out<=1;
   11616: out<=0;
   11617: out<=1;
   11618: out<=0;
   11619: out<=1;
   11620: out<=1;
   11621: out<=1;
   11622: out<=0;
   11623: out<=0;
   11624: out<=1;
   11625: out<=1;
   11626: out<=1;
   11627: out<=1;
   11628: out<=0;
   11629: out<=1;
   11630: out<=1;
   11631: out<=0;
   11632: out<=1;
   11633: out<=1;
   11634: out<=0;
   11635: out<=0;
   11636: out<=1;
   11637: out<=0;
   11638: out<=1;
   11639: out<=0;
   11640: out<=1;
   11641: out<=0;
   11642: out<=0;
   11643: out<=1;
   11644: out<=1;
   11645: out<=1;
   11646: out<=1;
   11647: out<=1;
   11648: out<=0;
   11649: out<=0;
   11650: out<=0;
   11651: out<=0;
   11652: out<=0;
   11653: out<=1;
   11654: out<=1;
   11655: out<=0;
   11656: out<=1;
   11657: out<=0;
   11658: out<=1;
   11659: out<=0;
   11660: out<=1;
   11661: out<=1;
   11662: out<=0;
   11663: out<=0;
   11664: out<=1;
   11665: out<=0;
   11666: out<=0;
   11667: out<=1;
   11668: out<=0;
   11669: out<=0;
   11670: out<=0;
   11671: out<=0;
   11672: out<=1;
   11673: out<=1;
   11674: out<=0;
   11675: out<=0;
   11676: out<=0;
   11677: out<=1;
   11678: out<=0;
   11679: out<=1;
   11680: out<=1;
   11681: out<=0;
   11682: out<=1;
   11683: out<=0;
   11684: out<=0;
   11685: out<=0;
   11686: out<=1;
   11687: out<=1;
   11688: out<=0;
   11689: out<=0;
   11690: out<=0;
   11691: out<=0;
   11692: out<=1;
   11693: out<=0;
   11694: out<=0;
   11695: out<=1;
   11696: out<=0;
   11697: out<=0;
   11698: out<=1;
   11699: out<=1;
   11700: out<=0;
   11701: out<=1;
   11702: out<=0;
   11703: out<=1;
   11704: out<=0;
   11705: out<=1;
   11706: out<=1;
   11707: out<=0;
   11708: out<=0;
   11709: out<=0;
   11710: out<=0;
   11711: out<=0;
   11712: out<=0;
   11713: out<=0;
   11714: out<=0;
   11715: out<=0;
   11716: out<=0;
   11717: out<=1;
   11718: out<=1;
   11719: out<=0;
   11720: out<=1;
   11721: out<=0;
   11722: out<=1;
   11723: out<=0;
   11724: out<=1;
   11725: out<=1;
   11726: out<=0;
   11727: out<=0;
   11728: out<=0;
   11729: out<=1;
   11730: out<=1;
   11731: out<=0;
   11732: out<=1;
   11733: out<=1;
   11734: out<=1;
   11735: out<=1;
   11736: out<=0;
   11737: out<=0;
   11738: out<=1;
   11739: out<=1;
   11740: out<=1;
   11741: out<=0;
   11742: out<=1;
   11743: out<=0;
   11744: out<=0;
   11745: out<=1;
   11746: out<=0;
   11747: out<=1;
   11748: out<=1;
   11749: out<=1;
   11750: out<=0;
   11751: out<=0;
   11752: out<=1;
   11753: out<=1;
   11754: out<=1;
   11755: out<=1;
   11756: out<=0;
   11757: out<=1;
   11758: out<=1;
   11759: out<=0;
   11760: out<=0;
   11761: out<=0;
   11762: out<=1;
   11763: out<=1;
   11764: out<=0;
   11765: out<=1;
   11766: out<=0;
   11767: out<=1;
   11768: out<=0;
   11769: out<=1;
   11770: out<=1;
   11771: out<=0;
   11772: out<=0;
   11773: out<=0;
   11774: out<=0;
   11775: out<=0;
   11776: out<=0;
   11777: out<=0;
   11778: out<=1;
   11779: out<=1;
   11780: out<=0;
   11781: out<=1;
   11782: out<=0;
   11783: out<=1;
   11784: out<=0;
   11785: out<=1;
   11786: out<=1;
   11787: out<=0;
   11788: out<=0;
   11789: out<=0;
   11790: out<=0;
   11791: out<=0;
   11792: out<=0;
   11793: out<=1;
   11794: out<=0;
   11795: out<=1;
   11796: out<=1;
   11797: out<=1;
   11798: out<=0;
   11799: out<=0;
   11800: out<=1;
   11801: out<=1;
   11802: out<=1;
   11803: out<=1;
   11804: out<=0;
   11805: out<=1;
   11806: out<=1;
   11807: out<=0;
   11808: out<=0;
   11809: out<=1;
   11810: out<=1;
   11811: out<=0;
   11812: out<=1;
   11813: out<=1;
   11814: out<=1;
   11815: out<=1;
   11816: out<=0;
   11817: out<=0;
   11818: out<=1;
   11819: out<=1;
   11820: out<=1;
   11821: out<=0;
   11822: out<=1;
   11823: out<=0;
   11824: out<=0;
   11825: out<=0;
   11826: out<=0;
   11827: out<=0;
   11828: out<=0;
   11829: out<=1;
   11830: out<=1;
   11831: out<=0;
   11832: out<=1;
   11833: out<=0;
   11834: out<=1;
   11835: out<=0;
   11836: out<=1;
   11837: out<=1;
   11838: out<=0;
   11839: out<=0;
   11840: out<=0;
   11841: out<=0;
   11842: out<=1;
   11843: out<=1;
   11844: out<=0;
   11845: out<=1;
   11846: out<=0;
   11847: out<=1;
   11848: out<=0;
   11849: out<=1;
   11850: out<=1;
   11851: out<=0;
   11852: out<=0;
   11853: out<=0;
   11854: out<=0;
   11855: out<=0;
   11856: out<=1;
   11857: out<=0;
   11858: out<=1;
   11859: out<=0;
   11860: out<=0;
   11861: out<=0;
   11862: out<=1;
   11863: out<=1;
   11864: out<=0;
   11865: out<=0;
   11866: out<=0;
   11867: out<=0;
   11868: out<=1;
   11869: out<=0;
   11870: out<=0;
   11871: out<=1;
   11872: out<=1;
   11873: out<=0;
   11874: out<=0;
   11875: out<=1;
   11876: out<=0;
   11877: out<=0;
   11878: out<=0;
   11879: out<=0;
   11880: out<=1;
   11881: out<=1;
   11882: out<=0;
   11883: out<=0;
   11884: out<=0;
   11885: out<=1;
   11886: out<=0;
   11887: out<=1;
   11888: out<=0;
   11889: out<=0;
   11890: out<=0;
   11891: out<=0;
   11892: out<=0;
   11893: out<=1;
   11894: out<=1;
   11895: out<=0;
   11896: out<=1;
   11897: out<=0;
   11898: out<=1;
   11899: out<=0;
   11900: out<=1;
   11901: out<=1;
   11902: out<=0;
   11903: out<=0;
   11904: out<=1;
   11905: out<=1;
   11906: out<=0;
   11907: out<=0;
   11908: out<=1;
   11909: out<=0;
   11910: out<=1;
   11911: out<=0;
   11912: out<=1;
   11913: out<=0;
   11914: out<=0;
   11915: out<=1;
   11916: out<=1;
   11917: out<=1;
   11918: out<=1;
   11919: out<=1;
   11920: out<=0;
   11921: out<=1;
   11922: out<=0;
   11923: out<=1;
   11924: out<=1;
   11925: out<=1;
   11926: out<=0;
   11927: out<=0;
   11928: out<=1;
   11929: out<=1;
   11930: out<=1;
   11931: out<=1;
   11932: out<=0;
   11933: out<=1;
   11934: out<=1;
   11935: out<=0;
   11936: out<=1;
   11937: out<=0;
   11938: out<=0;
   11939: out<=1;
   11940: out<=0;
   11941: out<=0;
   11942: out<=0;
   11943: out<=0;
   11944: out<=1;
   11945: out<=1;
   11946: out<=0;
   11947: out<=0;
   11948: out<=0;
   11949: out<=1;
   11950: out<=0;
   11951: out<=1;
   11952: out<=0;
   11953: out<=0;
   11954: out<=0;
   11955: out<=0;
   11956: out<=0;
   11957: out<=1;
   11958: out<=1;
   11959: out<=0;
   11960: out<=1;
   11961: out<=0;
   11962: out<=1;
   11963: out<=0;
   11964: out<=1;
   11965: out<=1;
   11966: out<=0;
   11967: out<=0;
   11968: out<=1;
   11969: out<=1;
   11970: out<=0;
   11971: out<=0;
   11972: out<=1;
   11973: out<=0;
   11974: out<=1;
   11975: out<=0;
   11976: out<=1;
   11977: out<=0;
   11978: out<=0;
   11979: out<=1;
   11980: out<=1;
   11981: out<=1;
   11982: out<=1;
   11983: out<=1;
   11984: out<=1;
   11985: out<=0;
   11986: out<=1;
   11987: out<=0;
   11988: out<=0;
   11989: out<=0;
   11990: out<=1;
   11991: out<=1;
   11992: out<=0;
   11993: out<=0;
   11994: out<=0;
   11995: out<=0;
   11996: out<=1;
   11997: out<=0;
   11998: out<=0;
   11999: out<=1;
   12000: out<=0;
   12001: out<=1;
   12002: out<=1;
   12003: out<=0;
   12004: out<=1;
   12005: out<=1;
   12006: out<=1;
   12007: out<=1;
   12008: out<=0;
   12009: out<=0;
   12010: out<=1;
   12011: out<=1;
   12012: out<=1;
   12013: out<=0;
   12014: out<=1;
   12015: out<=0;
   12016: out<=0;
   12017: out<=0;
   12018: out<=0;
   12019: out<=0;
   12020: out<=0;
   12021: out<=1;
   12022: out<=1;
   12023: out<=0;
   12024: out<=1;
   12025: out<=0;
   12026: out<=1;
   12027: out<=0;
   12028: out<=1;
   12029: out<=1;
   12030: out<=0;
   12031: out<=0;
   12032: out<=1;
   12033: out<=0;
   12034: out<=1;
   12035: out<=0;
   12036: out<=0;
   12037: out<=0;
   12038: out<=1;
   12039: out<=1;
   12040: out<=0;
   12041: out<=0;
   12042: out<=0;
   12043: out<=0;
   12044: out<=1;
   12045: out<=0;
   12046: out<=0;
   12047: out<=1;
   12048: out<=0;
   12049: out<=0;
   12050: out<=1;
   12051: out<=1;
   12052: out<=0;
   12053: out<=1;
   12054: out<=0;
   12055: out<=1;
   12056: out<=0;
   12057: out<=1;
   12058: out<=1;
   12059: out<=0;
   12060: out<=0;
   12061: out<=0;
   12062: out<=0;
   12063: out<=0;
   12064: out<=0;
   12065: out<=0;
   12066: out<=0;
   12067: out<=0;
   12068: out<=0;
   12069: out<=1;
   12070: out<=1;
   12071: out<=0;
   12072: out<=1;
   12073: out<=0;
   12074: out<=1;
   12075: out<=0;
   12076: out<=1;
   12077: out<=1;
   12078: out<=0;
   12079: out<=0;
   12080: out<=1;
   12081: out<=0;
   12082: out<=0;
   12083: out<=1;
   12084: out<=0;
   12085: out<=0;
   12086: out<=0;
   12087: out<=0;
   12088: out<=1;
   12089: out<=1;
   12090: out<=0;
   12091: out<=0;
   12092: out<=0;
   12093: out<=1;
   12094: out<=0;
   12095: out<=1;
   12096: out<=0;
   12097: out<=1;
   12098: out<=0;
   12099: out<=1;
   12100: out<=1;
   12101: out<=1;
   12102: out<=0;
   12103: out<=0;
   12104: out<=1;
   12105: out<=1;
   12106: out<=1;
   12107: out<=1;
   12108: out<=0;
   12109: out<=1;
   12110: out<=1;
   12111: out<=0;
   12112: out<=0;
   12113: out<=0;
   12114: out<=1;
   12115: out<=1;
   12116: out<=0;
   12117: out<=1;
   12118: out<=0;
   12119: out<=1;
   12120: out<=0;
   12121: out<=1;
   12122: out<=1;
   12123: out<=0;
   12124: out<=0;
   12125: out<=0;
   12126: out<=0;
   12127: out<=0;
   12128: out<=0;
   12129: out<=0;
   12130: out<=0;
   12131: out<=0;
   12132: out<=0;
   12133: out<=1;
   12134: out<=1;
   12135: out<=0;
   12136: out<=1;
   12137: out<=0;
   12138: out<=1;
   12139: out<=0;
   12140: out<=1;
   12141: out<=1;
   12142: out<=0;
   12143: out<=0;
   12144: out<=0;
   12145: out<=1;
   12146: out<=1;
   12147: out<=0;
   12148: out<=1;
   12149: out<=1;
   12150: out<=1;
   12151: out<=1;
   12152: out<=0;
   12153: out<=0;
   12154: out<=1;
   12155: out<=1;
   12156: out<=1;
   12157: out<=0;
   12158: out<=1;
   12159: out<=0;
   12160: out<=1;
   12161: out<=0;
   12162: out<=1;
   12163: out<=0;
   12164: out<=0;
   12165: out<=0;
   12166: out<=1;
   12167: out<=1;
   12168: out<=0;
   12169: out<=0;
   12170: out<=0;
   12171: out<=0;
   12172: out<=1;
   12173: out<=0;
   12174: out<=0;
   12175: out<=1;
   12176: out<=1;
   12177: out<=1;
   12178: out<=0;
   12179: out<=0;
   12180: out<=1;
   12181: out<=0;
   12182: out<=1;
   12183: out<=0;
   12184: out<=1;
   12185: out<=0;
   12186: out<=0;
   12187: out<=1;
   12188: out<=1;
   12189: out<=1;
   12190: out<=1;
   12191: out<=1;
   12192: out<=0;
   12193: out<=0;
   12194: out<=0;
   12195: out<=0;
   12196: out<=0;
   12197: out<=1;
   12198: out<=1;
   12199: out<=0;
   12200: out<=1;
   12201: out<=0;
   12202: out<=1;
   12203: out<=0;
   12204: out<=1;
   12205: out<=1;
   12206: out<=0;
   12207: out<=0;
   12208: out<=0;
   12209: out<=1;
   12210: out<=1;
   12211: out<=0;
   12212: out<=1;
   12213: out<=1;
   12214: out<=1;
   12215: out<=1;
   12216: out<=0;
   12217: out<=0;
   12218: out<=1;
   12219: out<=1;
   12220: out<=1;
   12221: out<=0;
   12222: out<=1;
   12223: out<=0;
   12224: out<=0;
   12225: out<=1;
   12226: out<=0;
   12227: out<=1;
   12228: out<=1;
   12229: out<=1;
   12230: out<=0;
   12231: out<=0;
   12232: out<=1;
   12233: out<=1;
   12234: out<=1;
   12235: out<=1;
   12236: out<=0;
   12237: out<=1;
   12238: out<=1;
   12239: out<=0;
   12240: out<=1;
   12241: out<=1;
   12242: out<=0;
   12243: out<=0;
   12244: out<=1;
   12245: out<=0;
   12246: out<=1;
   12247: out<=0;
   12248: out<=1;
   12249: out<=0;
   12250: out<=0;
   12251: out<=1;
   12252: out<=1;
   12253: out<=1;
   12254: out<=1;
   12255: out<=1;
   12256: out<=0;
   12257: out<=0;
   12258: out<=0;
   12259: out<=0;
   12260: out<=0;
   12261: out<=1;
   12262: out<=1;
   12263: out<=0;
   12264: out<=1;
   12265: out<=0;
   12266: out<=1;
   12267: out<=0;
   12268: out<=1;
   12269: out<=1;
   12270: out<=0;
   12271: out<=0;
   12272: out<=1;
   12273: out<=0;
   12274: out<=0;
   12275: out<=1;
   12276: out<=0;
   12277: out<=0;
   12278: out<=0;
   12279: out<=0;
   12280: out<=1;
   12281: out<=1;
   12282: out<=0;
   12283: out<=0;
   12284: out<=0;
   12285: out<=1;
   12286: out<=0;
   12287: out<=1;
   12288: out<=1;
   12289: out<=0;
   12290: out<=1;
   12291: out<=0;
   12292: out<=1;
   12293: out<=1;
   12294: out<=0;
   12295: out<=0;
   12296: out<=0;
   12297: out<=0;
   12298: out<=0;
   12299: out<=0;
   12300: out<=0;
   12301: out<=1;
   12302: out<=1;
   12303: out<=0;
   12304: out<=0;
   12305: out<=0;
   12306: out<=1;
   12307: out<=1;
   12308: out<=1;
   12309: out<=0;
   12310: out<=1;
   12311: out<=0;
   12312: out<=0;
   12313: out<=1;
   12314: out<=1;
   12315: out<=0;
   12316: out<=1;
   12317: out<=1;
   12318: out<=1;
   12319: out<=1;
   12320: out<=1;
   12321: out<=1;
   12322: out<=1;
   12323: out<=1;
   12324: out<=0;
   12325: out<=1;
   12326: out<=1;
   12327: out<=0;
   12328: out<=0;
   12329: out<=1;
   12330: out<=0;
   12331: out<=1;
   12332: out<=1;
   12333: out<=1;
   12334: out<=0;
   12335: out<=0;
   12336: out<=0;
   12337: out<=1;
   12338: out<=1;
   12339: out<=0;
   12340: out<=0;
   12341: out<=0;
   12342: out<=0;
   12343: out<=0;
   12344: out<=0;
   12345: out<=0;
   12346: out<=1;
   12347: out<=1;
   12348: out<=0;
   12349: out<=1;
   12350: out<=0;
   12351: out<=1;
   12352: out<=0;
   12353: out<=1;
   12354: out<=0;
   12355: out<=1;
   12356: out<=0;
   12357: out<=0;
   12358: out<=1;
   12359: out<=1;
   12360: out<=1;
   12361: out<=1;
   12362: out<=1;
   12363: out<=1;
   12364: out<=1;
   12365: out<=0;
   12366: out<=0;
   12367: out<=1;
   12368: out<=0;
   12369: out<=0;
   12370: out<=1;
   12371: out<=1;
   12372: out<=1;
   12373: out<=0;
   12374: out<=1;
   12375: out<=0;
   12376: out<=0;
   12377: out<=1;
   12378: out<=1;
   12379: out<=0;
   12380: out<=1;
   12381: out<=1;
   12382: out<=1;
   12383: out<=1;
   12384: out<=1;
   12385: out<=1;
   12386: out<=1;
   12387: out<=1;
   12388: out<=0;
   12389: out<=1;
   12390: out<=1;
   12391: out<=0;
   12392: out<=0;
   12393: out<=1;
   12394: out<=0;
   12395: out<=1;
   12396: out<=1;
   12397: out<=1;
   12398: out<=0;
   12399: out<=0;
   12400: out<=1;
   12401: out<=0;
   12402: out<=0;
   12403: out<=1;
   12404: out<=1;
   12405: out<=1;
   12406: out<=1;
   12407: out<=1;
   12408: out<=1;
   12409: out<=1;
   12410: out<=0;
   12411: out<=0;
   12412: out<=1;
   12413: out<=0;
   12414: out<=1;
   12415: out<=0;
   12416: out<=1;
   12417: out<=0;
   12418: out<=1;
   12419: out<=0;
   12420: out<=1;
   12421: out<=1;
   12422: out<=0;
   12423: out<=0;
   12424: out<=0;
   12425: out<=0;
   12426: out<=0;
   12427: out<=0;
   12428: out<=0;
   12429: out<=1;
   12430: out<=1;
   12431: out<=0;
   12432: out<=1;
   12433: out<=1;
   12434: out<=0;
   12435: out<=0;
   12436: out<=0;
   12437: out<=1;
   12438: out<=0;
   12439: out<=1;
   12440: out<=1;
   12441: out<=0;
   12442: out<=0;
   12443: out<=1;
   12444: out<=0;
   12445: out<=0;
   12446: out<=0;
   12447: out<=0;
   12448: out<=1;
   12449: out<=1;
   12450: out<=1;
   12451: out<=1;
   12452: out<=0;
   12453: out<=1;
   12454: out<=1;
   12455: out<=0;
   12456: out<=0;
   12457: out<=1;
   12458: out<=0;
   12459: out<=1;
   12460: out<=1;
   12461: out<=1;
   12462: out<=0;
   12463: out<=0;
   12464: out<=1;
   12465: out<=0;
   12466: out<=0;
   12467: out<=1;
   12468: out<=1;
   12469: out<=1;
   12470: out<=1;
   12471: out<=1;
   12472: out<=1;
   12473: out<=1;
   12474: out<=0;
   12475: out<=0;
   12476: out<=1;
   12477: out<=0;
   12478: out<=1;
   12479: out<=0;
   12480: out<=0;
   12481: out<=1;
   12482: out<=0;
   12483: out<=1;
   12484: out<=0;
   12485: out<=0;
   12486: out<=1;
   12487: out<=1;
   12488: out<=1;
   12489: out<=1;
   12490: out<=1;
   12491: out<=1;
   12492: out<=1;
   12493: out<=0;
   12494: out<=0;
   12495: out<=1;
   12496: out<=1;
   12497: out<=1;
   12498: out<=0;
   12499: out<=0;
   12500: out<=0;
   12501: out<=1;
   12502: out<=0;
   12503: out<=1;
   12504: out<=1;
   12505: out<=0;
   12506: out<=0;
   12507: out<=1;
   12508: out<=0;
   12509: out<=0;
   12510: out<=0;
   12511: out<=0;
   12512: out<=1;
   12513: out<=1;
   12514: out<=1;
   12515: out<=1;
   12516: out<=0;
   12517: out<=1;
   12518: out<=1;
   12519: out<=0;
   12520: out<=0;
   12521: out<=1;
   12522: out<=0;
   12523: out<=1;
   12524: out<=1;
   12525: out<=1;
   12526: out<=0;
   12527: out<=0;
   12528: out<=0;
   12529: out<=1;
   12530: out<=1;
   12531: out<=0;
   12532: out<=0;
   12533: out<=0;
   12534: out<=0;
   12535: out<=0;
   12536: out<=0;
   12537: out<=0;
   12538: out<=1;
   12539: out<=1;
   12540: out<=0;
   12541: out<=1;
   12542: out<=0;
   12543: out<=1;
   12544: out<=0;
   12545: out<=0;
   12546: out<=1;
   12547: out<=1;
   12548: out<=1;
   12549: out<=0;
   12550: out<=1;
   12551: out<=0;
   12552: out<=0;
   12553: out<=1;
   12554: out<=1;
   12555: out<=0;
   12556: out<=1;
   12557: out<=1;
   12558: out<=1;
   12559: out<=1;
   12560: out<=0;
   12561: out<=1;
   12562: out<=0;
   12563: out<=1;
   12564: out<=0;
   12565: out<=0;
   12566: out<=1;
   12567: out<=1;
   12568: out<=1;
   12569: out<=1;
   12570: out<=1;
   12571: out<=1;
   12572: out<=1;
   12573: out<=0;
   12574: out<=0;
   12575: out<=1;
   12576: out<=1;
   12577: out<=0;
   12578: out<=0;
   12579: out<=1;
   12580: out<=1;
   12581: out<=1;
   12582: out<=1;
   12583: out<=1;
   12584: out<=1;
   12585: out<=1;
   12586: out<=0;
   12587: out<=0;
   12588: out<=1;
   12589: out<=0;
   12590: out<=1;
   12591: out<=0;
   12592: out<=1;
   12593: out<=1;
   12594: out<=1;
   12595: out<=1;
   12596: out<=0;
   12597: out<=1;
   12598: out<=1;
   12599: out<=0;
   12600: out<=0;
   12601: out<=1;
   12602: out<=0;
   12603: out<=1;
   12604: out<=1;
   12605: out<=1;
   12606: out<=0;
   12607: out<=0;
   12608: out<=0;
   12609: out<=0;
   12610: out<=1;
   12611: out<=1;
   12612: out<=1;
   12613: out<=0;
   12614: out<=1;
   12615: out<=0;
   12616: out<=0;
   12617: out<=1;
   12618: out<=1;
   12619: out<=0;
   12620: out<=1;
   12621: out<=1;
   12622: out<=1;
   12623: out<=1;
   12624: out<=1;
   12625: out<=0;
   12626: out<=1;
   12627: out<=0;
   12628: out<=1;
   12629: out<=1;
   12630: out<=0;
   12631: out<=0;
   12632: out<=0;
   12633: out<=0;
   12634: out<=0;
   12635: out<=0;
   12636: out<=0;
   12637: out<=1;
   12638: out<=1;
   12639: out<=0;
   12640: out<=0;
   12641: out<=1;
   12642: out<=1;
   12643: out<=0;
   12644: out<=0;
   12645: out<=0;
   12646: out<=0;
   12647: out<=0;
   12648: out<=0;
   12649: out<=0;
   12650: out<=1;
   12651: out<=1;
   12652: out<=0;
   12653: out<=1;
   12654: out<=0;
   12655: out<=1;
   12656: out<=1;
   12657: out<=1;
   12658: out<=1;
   12659: out<=1;
   12660: out<=0;
   12661: out<=1;
   12662: out<=1;
   12663: out<=0;
   12664: out<=0;
   12665: out<=1;
   12666: out<=0;
   12667: out<=1;
   12668: out<=1;
   12669: out<=1;
   12670: out<=0;
   12671: out<=0;
   12672: out<=1;
   12673: out<=1;
   12674: out<=0;
   12675: out<=0;
   12676: out<=0;
   12677: out<=1;
   12678: out<=0;
   12679: out<=1;
   12680: out<=1;
   12681: out<=0;
   12682: out<=0;
   12683: out<=1;
   12684: out<=0;
   12685: out<=0;
   12686: out<=0;
   12687: out<=0;
   12688: out<=0;
   12689: out<=1;
   12690: out<=0;
   12691: out<=1;
   12692: out<=0;
   12693: out<=0;
   12694: out<=1;
   12695: out<=1;
   12696: out<=1;
   12697: out<=1;
   12698: out<=1;
   12699: out<=1;
   12700: out<=1;
   12701: out<=0;
   12702: out<=0;
   12703: out<=1;
   12704: out<=0;
   12705: out<=1;
   12706: out<=1;
   12707: out<=0;
   12708: out<=0;
   12709: out<=0;
   12710: out<=0;
   12711: out<=0;
   12712: out<=0;
   12713: out<=0;
   12714: out<=1;
   12715: out<=1;
   12716: out<=0;
   12717: out<=1;
   12718: out<=0;
   12719: out<=1;
   12720: out<=1;
   12721: out<=1;
   12722: out<=1;
   12723: out<=1;
   12724: out<=0;
   12725: out<=1;
   12726: out<=1;
   12727: out<=0;
   12728: out<=0;
   12729: out<=1;
   12730: out<=0;
   12731: out<=1;
   12732: out<=1;
   12733: out<=1;
   12734: out<=0;
   12735: out<=0;
   12736: out<=1;
   12737: out<=1;
   12738: out<=0;
   12739: out<=0;
   12740: out<=0;
   12741: out<=1;
   12742: out<=0;
   12743: out<=1;
   12744: out<=1;
   12745: out<=0;
   12746: out<=0;
   12747: out<=1;
   12748: out<=0;
   12749: out<=0;
   12750: out<=0;
   12751: out<=0;
   12752: out<=1;
   12753: out<=0;
   12754: out<=1;
   12755: out<=0;
   12756: out<=1;
   12757: out<=1;
   12758: out<=0;
   12759: out<=0;
   12760: out<=0;
   12761: out<=0;
   12762: out<=0;
   12763: out<=0;
   12764: out<=0;
   12765: out<=1;
   12766: out<=1;
   12767: out<=0;
   12768: out<=1;
   12769: out<=0;
   12770: out<=0;
   12771: out<=1;
   12772: out<=1;
   12773: out<=1;
   12774: out<=1;
   12775: out<=1;
   12776: out<=1;
   12777: out<=1;
   12778: out<=0;
   12779: out<=0;
   12780: out<=1;
   12781: out<=0;
   12782: out<=1;
   12783: out<=0;
   12784: out<=1;
   12785: out<=1;
   12786: out<=1;
   12787: out<=1;
   12788: out<=0;
   12789: out<=1;
   12790: out<=1;
   12791: out<=0;
   12792: out<=0;
   12793: out<=1;
   12794: out<=0;
   12795: out<=1;
   12796: out<=1;
   12797: out<=1;
   12798: out<=0;
   12799: out<=0;
   12800: out<=1;
   12801: out<=1;
   12802: out<=1;
   12803: out<=1;
   12804: out<=0;
   12805: out<=1;
   12806: out<=1;
   12807: out<=0;
   12808: out<=0;
   12809: out<=1;
   12810: out<=0;
   12811: out<=1;
   12812: out<=1;
   12813: out<=1;
   12814: out<=0;
   12815: out<=0;
   12816: out<=1;
   12817: out<=0;
   12818: out<=0;
   12819: out<=1;
   12820: out<=1;
   12821: out<=1;
   12822: out<=1;
   12823: out<=1;
   12824: out<=1;
   12825: out<=1;
   12826: out<=0;
   12827: out<=0;
   12828: out<=1;
   12829: out<=0;
   12830: out<=1;
   12831: out<=0;
   12832: out<=1;
   12833: out<=0;
   12834: out<=1;
   12835: out<=0;
   12836: out<=1;
   12837: out<=1;
   12838: out<=0;
   12839: out<=0;
   12840: out<=0;
   12841: out<=0;
   12842: out<=0;
   12843: out<=0;
   12844: out<=0;
   12845: out<=1;
   12846: out<=1;
   12847: out<=0;
   12848: out<=1;
   12849: out<=1;
   12850: out<=0;
   12851: out<=0;
   12852: out<=0;
   12853: out<=1;
   12854: out<=0;
   12855: out<=1;
   12856: out<=1;
   12857: out<=0;
   12858: out<=0;
   12859: out<=1;
   12860: out<=0;
   12861: out<=0;
   12862: out<=0;
   12863: out<=0;
   12864: out<=1;
   12865: out<=1;
   12866: out<=1;
   12867: out<=1;
   12868: out<=0;
   12869: out<=1;
   12870: out<=1;
   12871: out<=0;
   12872: out<=0;
   12873: out<=1;
   12874: out<=0;
   12875: out<=1;
   12876: out<=1;
   12877: out<=1;
   12878: out<=0;
   12879: out<=0;
   12880: out<=0;
   12881: out<=1;
   12882: out<=1;
   12883: out<=0;
   12884: out<=0;
   12885: out<=0;
   12886: out<=0;
   12887: out<=0;
   12888: out<=0;
   12889: out<=0;
   12890: out<=1;
   12891: out<=1;
   12892: out<=0;
   12893: out<=1;
   12894: out<=0;
   12895: out<=1;
   12896: out<=0;
   12897: out<=1;
   12898: out<=0;
   12899: out<=1;
   12900: out<=0;
   12901: out<=0;
   12902: out<=1;
   12903: out<=1;
   12904: out<=1;
   12905: out<=1;
   12906: out<=1;
   12907: out<=1;
   12908: out<=1;
   12909: out<=0;
   12910: out<=0;
   12911: out<=1;
   12912: out<=1;
   12913: out<=1;
   12914: out<=0;
   12915: out<=0;
   12916: out<=0;
   12917: out<=1;
   12918: out<=0;
   12919: out<=1;
   12920: out<=1;
   12921: out<=0;
   12922: out<=0;
   12923: out<=1;
   12924: out<=0;
   12925: out<=0;
   12926: out<=0;
   12927: out<=0;
   12928: out<=1;
   12929: out<=1;
   12930: out<=1;
   12931: out<=1;
   12932: out<=0;
   12933: out<=1;
   12934: out<=1;
   12935: out<=0;
   12936: out<=0;
   12937: out<=1;
   12938: out<=0;
   12939: out<=1;
   12940: out<=1;
   12941: out<=1;
   12942: out<=0;
   12943: out<=0;
   12944: out<=0;
   12945: out<=1;
   12946: out<=1;
   12947: out<=0;
   12948: out<=0;
   12949: out<=0;
   12950: out<=0;
   12951: out<=0;
   12952: out<=0;
   12953: out<=0;
   12954: out<=1;
   12955: out<=1;
   12956: out<=0;
   12957: out<=1;
   12958: out<=0;
   12959: out<=1;
   12960: out<=1;
   12961: out<=0;
   12962: out<=1;
   12963: out<=0;
   12964: out<=1;
   12965: out<=1;
   12966: out<=0;
   12967: out<=0;
   12968: out<=0;
   12969: out<=0;
   12970: out<=0;
   12971: out<=0;
   12972: out<=0;
   12973: out<=1;
   12974: out<=1;
   12975: out<=0;
   12976: out<=0;
   12977: out<=0;
   12978: out<=1;
   12979: out<=1;
   12980: out<=1;
   12981: out<=0;
   12982: out<=1;
   12983: out<=0;
   12984: out<=0;
   12985: out<=1;
   12986: out<=1;
   12987: out<=0;
   12988: out<=1;
   12989: out<=1;
   12990: out<=1;
   12991: out<=1;
   12992: out<=1;
   12993: out<=1;
   12994: out<=1;
   12995: out<=1;
   12996: out<=0;
   12997: out<=1;
   12998: out<=1;
   12999: out<=0;
   13000: out<=0;
   13001: out<=1;
   13002: out<=0;
   13003: out<=1;
   13004: out<=1;
   13005: out<=1;
   13006: out<=0;
   13007: out<=0;
   13008: out<=1;
   13009: out<=0;
   13010: out<=0;
   13011: out<=1;
   13012: out<=1;
   13013: out<=1;
   13014: out<=1;
   13015: out<=1;
   13016: out<=1;
   13017: out<=1;
   13018: out<=0;
   13019: out<=0;
   13020: out<=1;
   13021: out<=0;
   13022: out<=1;
   13023: out<=0;
   13024: out<=0;
   13025: out<=1;
   13026: out<=0;
   13027: out<=1;
   13028: out<=0;
   13029: out<=0;
   13030: out<=1;
   13031: out<=1;
   13032: out<=1;
   13033: out<=1;
   13034: out<=1;
   13035: out<=1;
   13036: out<=1;
   13037: out<=0;
   13038: out<=0;
   13039: out<=1;
   13040: out<=0;
   13041: out<=0;
   13042: out<=1;
   13043: out<=1;
   13044: out<=1;
   13045: out<=0;
   13046: out<=1;
   13047: out<=0;
   13048: out<=0;
   13049: out<=1;
   13050: out<=1;
   13051: out<=0;
   13052: out<=1;
   13053: out<=1;
   13054: out<=1;
   13055: out<=1;
   13056: out<=0;
   13057: out<=1;
   13058: out<=1;
   13059: out<=0;
   13060: out<=0;
   13061: out<=0;
   13062: out<=0;
   13063: out<=0;
   13064: out<=0;
   13065: out<=0;
   13066: out<=1;
   13067: out<=1;
   13068: out<=0;
   13069: out<=1;
   13070: out<=0;
   13071: out<=1;
   13072: out<=1;
   13073: out<=1;
   13074: out<=1;
   13075: out<=1;
   13076: out<=0;
   13077: out<=1;
   13078: out<=1;
   13079: out<=0;
   13080: out<=0;
   13081: out<=1;
   13082: out<=0;
   13083: out<=1;
   13084: out<=1;
   13085: out<=1;
   13086: out<=0;
   13087: out<=0;
   13088: out<=1;
   13089: out<=1;
   13090: out<=0;
   13091: out<=0;
   13092: out<=0;
   13093: out<=1;
   13094: out<=0;
   13095: out<=1;
   13096: out<=1;
   13097: out<=0;
   13098: out<=0;
   13099: out<=1;
   13100: out<=0;
   13101: out<=0;
   13102: out<=0;
   13103: out<=0;
   13104: out<=0;
   13105: out<=1;
   13106: out<=0;
   13107: out<=1;
   13108: out<=0;
   13109: out<=0;
   13110: out<=1;
   13111: out<=1;
   13112: out<=1;
   13113: out<=1;
   13114: out<=1;
   13115: out<=1;
   13116: out<=1;
   13117: out<=0;
   13118: out<=0;
   13119: out<=1;
   13120: out<=1;
   13121: out<=0;
   13122: out<=0;
   13123: out<=1;
   13124: out<=1;
   13125: out<=1;
   13126: out<=1;
   13127: out<=1;
   13128: out<=1;
   13129: out<=1;
   13130: out<=0;
   13131: out<=0;
   13132: out<=1;
   13133: out<=0;
   13134: out<=1;
   13135: out<=0;
   13136: out<=1;
   13137: out<=1;
   13138: out<=1;
   13139: out<=1;
   13140: out<=0;
   13141: out<=1;
   13142: out<=1;
   13143: out<=0;
   13144: out<=0;
   13145: out<=1;
   13146: out<=0;
   13147: out<=1;
   13148: out<=1;
   13149: out<=1;
   13150: out<=0;
   13151: out<=0;
   13152: out<=1;
   13153: out<=1;
   13154: out<=0;
   13155: out<=0;
   13156: out<=0;
   13157: out<=1;
   13158: out<=0;
   13159: out<=1;
   13160: out<=1;
   13161: out<=0;
   13162: out<=0;
   13163: out<=1;
   13164: out<=0;
   13165: out<=0;
   13166: out<=0;
   13167: out<=0;
   13168: out<=1;
   13169: out<=0;
   13170: out<=1;
   13171: out<=0;
   13172: out<=1;
   13173: out<=1;
   13174: out<=0;
   13175: out<=0;
   13176: out<=0;
   13177: out<=0;
   13178: out<=0;
   13179: out<=0;
   13180: out<=0;
   13181: out<=1;
   13182: out<=1;
   13183: out<=0;
   13184: out<=1;
   13185: out<=0;
   13186: out<=0;
   13187: out<=1;
   13188: out<=1;
   13189: out<=1;
   13190: out<=1;
   13191: out<=1;
   13192: out<=1;
   13193: out<=1;
   13194: out<=0;
   13195: out<=0;
   13196: out<=1;
   13197: out<=0;
   13198: out<=1;
   13199: out<=0;
   13200: out<=1;
   13201: out<=1;
   13202: out<=1;
   13203: out<=1;
   13204: out<=0;
   13205: out<=1;
   13206: out<=1;
   13207: out<=0;
   13208: out<=0;
   13209: out<=1;
   13210: out<=0;
   13211: out<=1;
   13212: out<=1;
   13213: out<=1;
   13214: out<=0;
   13215: out<=0;
   13216: out<=0;
   13217: out<=0;
   13218: out<=1;
   13219: out<=1;
   13220: out<=1;
   13221: out<=0;
   13222: out<=1;
   13223: out<=0;
   13224: out<=0;
   13225: out<=1;
   13226: out<=1;
   13227: out<=0;
   13228: out<=1;
   13229: out<=1;
   13230: out<=1;
   13231: out<=1;
   13232: out<=0;
   13233: out<=1;
   13234: out<=0;
   13235: out<=1;
   13236: out<=0;
   13237: out<=0;
   13238: out<=1;
   13239: out<=1;
   13240: out<=1;
   13241: out<=1;
   13242: out<=1;
   13243: out<=1;
   13244: out<=1;
   13245: out<=0;
   13246: out<=0;
   13247: out<=1;
   13248: out<=0;
   13249: out<=1;
   13250: out<=1;
   13251: out<=0;
   13252: out<=0;
   13253: out<=0;
   13254: out<=0;
   13255: out<=0;
   13256: out<=0;
   13257: out<=0;
   13258: out<=1;
   13259: out<=1;
   13260: out<=0;
   13261: out<=1;
   13262: out<=0;
   13263: out<=1;
   13264: out<=1;
   13265: out<=1;
   13266: out<=1;
   13267: out<=1;
   13268: out<=0;
   13269: out<=1;
   13270: out<=1;
   13271: out<=0;
   13272: out<=0;
   13273: out<=1;
   13274: out<=0;
   13275: out<=1;
   13276: out<=1;
   13277: out<=1;
   13278: out<=0;
   13279: out<=0;
   13280: out<=0;
   13281: out<=0;
   13282: out<=1;
   13283: out<=1;
   13284: out<=1;
   13285: out<=0;
   13286: out<=1;
   13287: out<=0;
   13288: out<=0;
   13289: out<=1;
   13290: out<=1;
   13291: out<=0;
   13292: out<=1;
   13293: out<=1;
   13294: out<=1;
   13295: out<=1;
   13296: out<=1;
   13297: out<=0;
   13298: out<=1;
   13299: out<=0;
   13300: out<=1;
   13301: out<=1;
   13302: out<=0;
   13303: out<=0;
   13304: out<=0;
   13305: out<=0;
   13306: out<=0;
   13307: out<=0;
   13308: out<=0;
   13309: out<=1;
   13310: out<=1;
   13311: out<=0;
   13312: out<=0;
   13313: out<=0;
   13314: out<=1;
   13315: out<=1;
   13316: out<=0;
   13317: out<=1;
   13318: out<=0;
   13319: out<=1;
   13320: out<=1;
   13321: out<=0;
   13322: out<=0;
   13323: out<=1;
   13324: out<=1;
   13325: out<=1;
   13326: out<=1;
   13327: out<=1;
   13328: out<=1;
   13329: out<=0;
   13330: out<=1;
   13331: out<=0;
   13332: out<=0;
   13333: out<=0;
   13334: out<=1;
   13335: out<=1;
   13336: out<=1;
   13337: out<=1;
   13338: out<=1;
   13339: out<=1;
   13340: out<=0;
   13341: out<=1;
   13342: out<=1;
   13343: out<=0;
   13344: out<=0;
   13345: out<=1;
   13346: out<=1;
   13347: out<=0;
   13348: out<=1;
   13349: out<=1;
   13350: out<=1;
   13351: out<=1;
   13352: out<=1;
   13353: out<=1;
   13354: out<=0;
   13355: out<=0;
   13356: out<=0;
   13357: out<=1;
   13358: out<=0;
   13359: out<=1;
   13360: out<=1;
   13361: out<=1;
   13362: out<=1;
   13363: out<=1;
   13364: out<=1;
   13365: out<=0;
   13366: out<=0;
   13367: out<=1;
   13368: out<=1;
   13369: out<=0;
   13370: out<=1;
   13371: out<=0;
   13372: out<=1;
   13373: out<=1;
   13374: out<=0;
   13375: out<=0;
   13376: out<=0;
   13377: out<=0;
   13378: out<=1;
   13379: out<=1;
   13380: out<=0;
   13381: out<=1;
   13382: out<=0;
   13383: out<=1;
   13384: out<=1;
   13385: out<=0;
   13386: out<=0;
   13387: out<=1;
   13388: out<=1;
   13389: out<=1;
   13390: out<=1;
   13391: out<=1;
   13392: out<=0;
   13393: out<=1;
   13394: out<=0;
   13395: out<=1;
   13396: out<=1;
   13397: out<=1;
   13398: out<=0;
   13399: out<=0;
   13400: out<=0;
   13401: out<=0;
   13402: out<=0;
   13403: out<=0;
   13404: out<=1;
   13405: out<=0;
   13406: out<=0;
   13407: out<=1;
   13408: out<=1;
   13409: out<=0;
   13410: out<=0;
   13411: out<=1;
   13412: out<=0;
   13413: out<=0;
   13414: out<=0;
   13415: out<=0;
   13416: out<=0;
   13417: out<=0;
   13418: out<=1;
   13419: out<=1;
   13420: out<=1;
   13421: out<=0;
   13422: out<=1;
   13423: out<=0;
   13424: out<=1;
   13425: out<=1;
   13426: out<=1;
   13427: out<=1;
   13428: out<=1;
   13429: out<=0;
   13430: out<=0;
   13431: out<=1;
   13432: out<=1;
   13433: out<=0;
   13434: out<=1;
   13435: out<=0;
   13436: out<=1;
   13437: out<=1;
   13438: out<=0;
   13439: out<=0;
   13440: out<=1;
   13441: out<=1;
   13442: out<=0;
   13443: out<=0;
   13444: out<=1;
   13445: out<=0;
   13446: out<=1;
   13447: out<=0;
   13448: out<=0;
   13449: out<=1;
   13450: out<=1;
   13451: out<=0;
   13452: out<=0;
   13453: out<=0;
   13454: out<=0;
   13455: out<=0;
   13456: out<=1;
   13457: out<=0;
   13458: out<=1;
   13459: out<=0;
   13460: out<=0;
   13461: out<=0;
   13462: out<=1;
   13463: out<=1;
   13464: out<=1;
   13465: out<=1;
   13466: out<=1;
   13467: out<=1;
   13468: out<=0;
   13469: out<=1;
   13470: out<=1;
   13471: out<=0;
   13472: out<=1;
   13473: out<=0;
   13474: out<=0;
   13475: out<=1;
   13476: out<=0;
   13477: out<=0;
   13478: out<=0;
   13479: out<=0;
   13480: out<=0;
   13481: out<=0;
   13482: out<=1;
   13483: out<=1;
   13484: out<=1;
   13485: out<=0;
   13486: out<=1;
   13487: out<=0;
   13488: out<=1;
   13489: out<=1;
   13490: out<=1;
   13491: out<=1;
   13492: out<=1;
   13493: out<=0;
   13494: out<=0;
   13495: out<=1;
   13496: out<=1;
   13497: out<=0;
   13498: out<=1;
   13499: out<=0;
   13500: out<=1;
   13501: out<=1;
   13502: out<=0;
   13503: out<=0;
   13504: out<=1;
   13505: out<=1;
   13506: out<=0;
   13507: out<=0;
   13508: out<=1;
   13509: out<=0;
   13510: out<=1;
   13511: out<=0;
   13512: out<=0;
   13513: out<=1;
   13514: out<=1;
   13515: out<=0;
   13516: out<=0;
   13517: out<=0;
   13518: out<=0;
   13519: out<=0;
   13520: out<=0;
   13521: out<=1;
   13522: out<=0;
   13523: out<=1;
   13524: out<=1;
   13525: out<=1;
   13526: out<=0;
   13527: out<=0;
   13528: out<=0;
   13529: out<=0;
   13530: out<=0;
   13531: out<=0;
   13532: out<=1;
   13533: out<=0;
   13534: out<=0;
   13535: out<=1;
   13536: out<=0;
   13537: out<=1;
   13538: out<=1;
   13539: out<=0;
   13540: out<=1;
   13541: out<=1;
   13542: out<=1;
   13543: out<=1;
   13544: out<=1;
   13545: out<=1;
   13546: out<=0;
   13547: out<=0;
   13548: out<=0;
   13549: out<=1;
   13550: out<=0;
   13551: out<=1;
   13552: out<=1;
   13553: out<=1;
   13554: out<=1;
   13555: out<=1;
   13556: out<=1;
   13557: out<=0;
   13558: out<=0;
   13559: out<=1;
   13560: out<=1;
   13561: out<=0;
   13562: out<=1;
   13563: out<=0;
   13564: out<=1;
   13565: out<=1;
   13566: out<=0;
   13567: out<=0;
   13568: out<=0;
   13569: out<=1;
   13570: out<=0;
   13571: out<=1;
   13572: out<=1;
   13573: out<=1;
   13574: out<=0;
   13575: out<=0;
   13576: out<=0;
   13577: out<=0;
   13578: out<=0;
   13579: out<=0;
   13580: out<=1;
   13581: out<=0;
   13582: out<=0;
   13583: out<=1;
   13584: out<=0;
   13585: out<=0;
   13586: out<=1;
   13587: out<=1;
   13588: out<=0;
   13589: out<=1;
   13590: out<=0;
   13591: out<=1;
   13592: out<=1;
   13593: out<=0;
   13594: out<=0;
   13595: out<=1;
   13596: out<=1;
   13597: out<=1;
   13598: out<=1;
   13599: out<=1;
   13600: out<=1;
   13601: out<=1;
   13602: out<=1;
   13603: out<=1;
   13604: out<=1;
   13605: out<=0;
   13606: out<=0;
   13607: out<=1;
   13608: out<=1;
   13609: out<=0;
   13610: out<=1;
   13611: out<=0;
   13612: out<=1;
   13613: out<=1;
   13614: out<=0;
   13615: out<=0;
   13616: out<=1;
   13617: out<=0;
   13618: out<=0;
   13619: out<=1;
   13620: out<=0;
   13621: out<=0;
   13622: out<=0;
   13623: out<=0;
   13624: out<=0;
   13625: out<=0;
   13626: out<=1;
   13627: out<=1;
   13628: out<=1;
   13629: out<=0;
   13630: out<=1;
   13631: out<=0;
   13632: out<=1;
   13633: out<=0;
   13634: out<=1;
   13635: out<=0;
   13636: out<=0;
   13637: out<=0;
   13638: out<=1;
   13639: out<=1;
   13640: out<=1;
   13641: out<=1;
   13642: out<=1;
   13643: out<=1;
   13644: out<=0;
   13645: out<=1;
   13646: out<=1;
   13647: out<=0;
   13648: out<=0;
   13649: out<=0;
   13650: out<=1;
   13651: out<=1;
   13652: out<=0;
   13653: out<=1;
   13654: out<=0;
   13655: out<=1;
   13656: out<=1;
   13657: out<=0;
   13658: out<=0;
   13659: out<=1;
   13660: out<=1;
   13661: out<=1;
   13662: out<=1;
   13663: out<=1;
   13664: out<=1;
   13665: out<=1;
   13666: out<=1;
   13667: out<=1;
   13668: out<=1;
   13669: out<=0;
   13670: out<=0;
   13671: out<=1;
   13672: out<=1;
   13673: out<=0;
   13674: out<=1;
   13675: out<=0;
   13676: out<=1;
   13677: out<=1;
   13678: out<=0;
   13679: out<=0;
   13680: out<=0;
   13681: out<=1;
   13682: out<=1;
   13683: out<=0;
   13684: out<=1;
   13685: out<=1;
   13686: out<=1;
   13687: out<=1;
   13688: out<=1;
   13689: out<=1;
   13690: out<=0;
   13691: out<=0;
   13692: out<=0;
   13693: out<=1;
   13694: out<=0;
   13695: out<=1;
   13696: out<=0;
   13697: out<=1;
   13698: out<=0;
   13699: out<=1;
   13700: out<=1;
   13701: out<=1;
   13702: out<=0;
   13703: out<=0;
   13704: out<=0;
   13705: out<=0;
   13706: out<=0;
   13707: out<=0;
   13708: out<=1;
   13709: out<=0;
   13710: out<=0;
   13711: out<=1;
   13712: out<=1;
   13713: out<=1;
   13714: out<=0;
   13715: out<=0;
   13716: out<=1;
   13717: out<=0;
   13718: out<=1;
   13719: out<=0;
   13720: out<=0;
   13721: out<=1;
   13722: out<=1;
   13723: out<=0;
   13724: out<=0;
   13725: out<=0;
   13726: out<=0;
   13727: out<=0;
   13728: out<=1;
   13729: out<=1;
   13730: out<=1;
   13731: out<=1;
   13732: out<=1;
   13733: out<=0;
   13734: out<=0;
   13735: out<=1;
   13736: out<=1;
   13737: out<=0;
   13738: out<=1;
   13739: out<=0;
   13740: out<=1;
   13741: out<=1;
   13742: out<=0;
   13743: out<=0;
   13744: out<=0;
   13745: out<=1;
   13746: out<=1;
   13747: out<=0;
   13748: out<=1;
   13749: out<=1;
   13750: out<=1;
   13751: out<=1;
   13752: out<=1;
   13753: out<=1;
   13754: out<=0;
   13755: out<=0;
   13756: out<=0;
   13757: out<=1;
   13758: out<=0;
   13759: out<=1;
   13760: out<=1;
   13761: out<=0;
   13762: out<=1;
   13763: out<=0;
   13764: out<=0;
   13765: out<=0;
   13766: out<=1;
   13767: out<=1;
   13768: out<=1;
   13769: out<=1;
   13770: out<=1;
   13771: out<=1;
   13772: out<=0;
   13773: out<=1;
   13774: out<=1;
   13775: out<=0;
   13776: out<=1;
   13777: out<=1;
   13778: out<=0;
   13779: out<=0;
   13780: out<=1;
   13781: out<=0;
   13782: out<=1;
   13783: out<=0;
   13784: out<=0;
   13785: out<=1;
   13786: out<=1;
   13787: out<=0;
   13788: out<=0;
   13789: out<=0;
   13790: out<=0;
   13791: out<=0;
   13792: out<=1;
   13793: out<=1;
   13794: out<=1;
   13795: out<=1;
   13796: out<=1;
   13797: out<=0;
   13798: out<=0;
   13799: out<=1;
   13800: out<=1;
   13801: out<=0;
   13802: out<=1;
   13803: out<=0;
   13804: out<=1;
   13805: out<=1;
   13806: out<=0;
   13807: out<=0;
   13808: out<=1;
   13809: out<=0;
   13810: out<=0;
   13811: out<=1;
   13812: out<=0;
   13813: out<=0;
   13814: out<=0;
   13815: out<=0;
   13816: out<=0;
   13817: out<=0;
   13818: out<=1;
   13819: out<=1;
   13820: out<=1;
   13821: out<=0;
   13822: out<=1;
   13823: out<=0;
   13824: out<=1;
   13825: out<=0;
   13826: out<=0;
   13827: out<=1;
   13828: out<=0;
   13829: out<=0;
   13830: out<=0;
   13831: out<=0;
   13832: out<=0;
   13833: out<=0;
   13834: out<=1;
   13835: out<=1;
   13836: out<=1;
   13837: out<=0;
   13838: out<=1;
   13839: out<=0;
   13840: out<=1;
   13841: out<=1;
   13842: out<=1;
   13843: out<=1;
   13844: out<=1;
   13845: out<=0;
   13846: out<=0;
   13847: out<=1;
   13848: out<=1;
   13849: out<=0;
   13850: out<=1;
   13851: out<=0;
   13852: out<=1;
   13853: out<=1;
   13854: out<=0;
   13855: out<=0;
   13856: out<=1;
   13857: out<=1;
   13858: out<=0;
   13859: out<=0;
   13860: out<=1;
   13861: out<=0;
   13862: out<=1;
   13863: out<=0;
   13864: out<=0;
   13865: out<=1;
   13866: out<=1;
   13867: out<=0;
   13868: out<=0;
   13869: out<=0;
   13870: out<=0;
   13871: out<=0;
   13872: out<=1;
   13873: out<=0;
   13874: out<=1;
   13875: out<=0;
   13876: out<=0;
   13877: out<=0;
   13878: out<=1;
   13879: out<=1;
   13880: out<=1;
   13881: out<=1;
   13882: out<=1;
   13883: out<=1;
   13884: out<=0;
   13885: out<=1;
   13886: out<=1;
   13887: out<=0;
   13888: out<=0;
   13889: out<=1;
   13890: out<=1;
   13891: out<=0;
   13892: out<=1;
   13893: out<=1;
   13894: out<=1;
   13895: out<=1;
   13896: out<=1;
   13897: out<=1;
   13898: out<=0;
   13899: out<=0;
   13900: out<=0;
   13901: out<=1;
   13902: out<=0;
   13903: out<=1;
   13904: out<=1;
   13905: out<=1;
   13906: out<=1;
   13907: out<=1;
   13908: out<=1;
   13909: out<=0;
   13910: out<=0;
   13911: out<=1;
   13912: out<=1;
   13913: out<=0;
   13914: out<=1;
   13915: out<=0;
   13916: out<=1;
   13917: out<=1;
   13918: out<=0;
   13919: out<=0;
   13920: out<=1;
   13921: out<=1;
   13922: out<=0;
   13923: out<=0;
   13924: out<=1;
   13925: out<=0;
   13926: out<=1;
   13927: out<=0;
   13928: out<=0;
   13929: out<=1;
   13930: out<=1;
   13931: out<=0;
   13932: out<=0;
   13933: out<=0;
   13934: out<=0;
   13935: out<=0;
   13936: out<=0;
   13937: out<=1;
   13938: out<=0;
   13939: out<=1;
   13940: out<=1;
   13941: out<=1;
   13942: out<=0;
   13943: out<=0;
   13944: out<=0;
   13945: out<=0;
   13946: out<=0;
   13947: out<=0;
   13948: out<=1;
   13949: out<=0;
   13950: out<=0;
   13951: out<=1;
   13952: out<=0;
   13953: out<=1;
   13954: out<=1;
   13955: out<=0;
   13956: out<=1;
   13957: out<=1;
   13958: out<=1;
   13959: out<=1;
   13960: out<=1;
   13961: out<=1;
   13962: out<=0;
   13963: out<=0;
   13964: out<=0;
   13965: out<=1;
   13966: out<=0;
   13967: out<=1;
   13968: out<=1;
   13969: out<=1;
   13970: out<=1;
   13971: out<=1;
   13972: out<=1;
   13973: out<=0;
   13974: out<=0;
   13975: out<=1;
   13976: out<=1;
   13977: out<=0;
   13978: out<=1;
   13979: out<=0;
   13980: out<=1;
   13981: out<=1;
   13982: out<=0;
   13983: out<=0;
   13984: out<=0;
   13985: out<=0;
   13986: out<=1;
   13987: out<=1;
   13988: out<=0;
   13989: out<=1;
   13990: out<=0;
   13991: out<=1;
   13992: out<=1;
   13993: out<=0;
   13994: out<=0;
   13995: out<=1;
   13996: out<=1;
   13997: out<=1;
   13998: out<=1;
   13999: out<=1;
   14000: out<=1;
   14001: out<=0;
   14002: out<=1;
   14003: out<=0;
   14004: out<=0;
   14005: out<=0;
   14006: out<=1;
   14007: out<=1;
   14008: out<=1;
   14009: out<=1;
   14010: out<=1;
   14011: out<=1;
   14012: out<=0;
   14013: out<=1;
   14014: out<=1;
   14015: out<=0;
   14016: out<=1;
   14017: out<=0;
   14018: out<=0;
   14019: out<=1;
   14020: out<=0;
   14021: out<=0;
   14022: out<=0;
   14023: out<=0;
   14024: out<=0;
   14025: out<=0;
   14026: out<=1;
   14027: out<=1;
   14028: out<=1;
   14029: out<=0;
   14030: out<=1;
   14031: out<=0;
   14032: out<=1;
   14033: out<=1;
   14034: out<=1;
   14035: out<=1;
   14036: out<=1;
   14037: out<=0;
   14038: out<=0;
   14039: out<=1;
   14040: out<=1;
   14041: out<=0;
   14042: out<=1;
   14043: out<=0;
   14044: out<=1;
   14045: out<=1;
   14046: out<=0;
   14047: out<=0;
   14048: out<=0;
   14049: out<=0;
   14050: out<=1;
   14051: out<=1;
   14052: out<=0;
   14053: out<=1;
   14054: out<=0;
   14055: out<=1;
   14056: out<=1;
   14057: out<=0;
   14058: out<=0;
   14059: out<=1;
   14060: out<=1;
   14061: out<=1;
   14062: out<=1;
   14063: out<=1;
   14064: out<=0;
   14065: out<=1;
   14066: out<=0;
   14067: out<=1;
   14068: out<=1;
   14069: out<=1;
   14070: out<=0;
   14071: out<=0;
   14072: out<=0;
   14073: out<=0;
   14074: out<=0;
   14075: out<=0;
   14076: out<=1;
   14077: out<=0;
   14078: out<=0;
   14079: out<=1;
   14080: out<=1;
   14081: out<=1;
   14082: out<=1;
   14083: out<=1;
   14084: out<=1;
   14085: out<=0;
   14086: out<=0;
   14087: out<=1;
   14088: out<=1;
   14089: out<=0;
   14090: out<=1;
   14091: out<=0;
   14092: out<=1;
   14093: out<=1;
   14094: out<=0;
   14095: out<=0;
   14096: out<=0;
   14097: out<=1;
   14098: out<=1;
   14099: out<=0;
   14100: out<=1;
   14101: out<=1;
   14102: out<=1;
   14103: out<=1;
   14104: out<=1;
   14105: out<=1;
   14106: out<=0;
   14107: out<=0;
   14108: out<=0;
   14109: out<=1;
   14110: out<=0;
   14111: out<=1;
   14112: out<=0;
   14113: out<=1;
   14114: out<=0;
   14115: out<=1;
   14116: out<=1;
   14117: out<=1;
   14118: out<=0;
   14119: out<=0;
   14120: out<=0;
   14121: out<=0;
   14122: out<=0;
   14123: out<=0;
   14124: out<=1;
   14125: out<=0;
   14126: out<=0;
   14127: out<=1;
   14128: out<=1;
   14129: out<=1;
   14130: out<=0;
   14131: out<=0;
   14132: out<=1;
   14133: out<=0;
   14134: out<=1;
   14135: out<=0;
   14136: out<=0;
   14137: out<=1;
   14138: out<=1;
   14139: out<=0;
   14140: out<=0;
   14141: out<=0;
   14142: out<=0;
   14143: out<=0;
   14144: out<=1;
   14145: out<=1;
   14146: out<=1;
   14147: out<=1;
   14148: out<=1;
   14149: out<=0;
   14150: out<=0;
   14151: out<=1;
   14152: out<=1;
   14153: out<=0;
   14154: out<=1;
   14155: out<=0;
   14156: out<=1;
   14157: out<=1;
   14158: out<=0;
   14159: out<=0;
   14160: out<=1;
   14161: out<=0;
   14162: out<=0;
   14163: out<=1;
   14164: out<=0;
   14165: out<=0;
   14166: out<=0;
   14167: out<=0;
   14168: out<=0;
   14169: out<=0;
   14170: out<=1;
   14171: out<=1;
   14172: out<=1;
   14173: out<=0;
   14174: out<=1;
   14175: out<=0;
   14176: out<=1;
   14177: out<=0;
   14178: out<=1;
   14179: out<=0;
   14180: out<=0;
   14181: out<=0;
   14182: out<=1;
   14183: out<=1;
   14184: out<=1;
   14185: out<=1;
   14186: out<=1;
   14187: out<=1;
   14188: out<=0;
   14189: out<=1;
   14190: out<=1;
   14191: out<=0;
   14192: out<=1;
   14193: out<=1;
   14194: out<=0;
   14195: out<=0;
   14196: out<=1;
   14197: out<=0;
   14198: out<=1;
   14199: out<=0;
   14200: out<=0;
   14201: out<=1;
   14202: out<=1;
   14203: out<=0;
   14204: out<=0;
   14205: out<=0;
   14206: out<=0;
   14207: out<=0;
   14208: out<=1;
   14209: out<=1;
   14210: out<=1;
   14211: out<=1;
   14212: out<=1;
   14213: out<=0;
   14214: out<=0;
   14215: out<=1;
   14216: out<=1;
   14217: out<=0;
   14218: out<=1;
   14219: out<=0;
   14220: out<=1;
   14221: out<=1;
   14222: out<=0;
   14223: out<=0;
   14224: out<=1;
   14225: out<=0;
   14226: out<=0;
   14227: out<=1;
   14228: out<=0;
   14229: out<=0;
   14230: out<=0;
   14231: out<=0;
   14232: out<=0;
   14233: out<=0;
   14234: out<=1;
   14235: out<=1;
   14236: out<=1;
   14237: out<=0;
   14238: out<=1;
   14239: out<=0;
   14240: out<=0;
   14241: out<=1;
   14242: out<=0;
   14243: out<=1;
   14244: out<=1;
   14245: out<=1;
   14246: out<=0;
   14247: out<=0;
   14248: out<=0;
   14249: out<=0;
   14250: out<=0;
   14251: out<=0;
   14252: out<=1;
   14253: out<=0;
   14254: out<=0;
   14255: out<=1;
   14256: out<=0;
   14257: out<=0;
   14258: out<=1;
   14259: out<=1;
   14260: out<=0;
   14261: out<=1;
   14262: out<=0;
   14263: out<=1;
   14264: out<=1;
   14265: out<=0;
   14266: out<=0;
   14267: out<=1;
   14268: out<=1;
   14269: out<=1;
   14270: out<=1;
   14271: out<=1;
   14272: out<=1;
   14273: out<=1;
   14274: out<=1;
   14275: out<=1;
   14276: out<=1;
   14277: out<=0;
   14278: out<=0;
   14279: out<=1;
   14280: out<=1;
   14281: out<=0;
   14282: out<=1;
   14283: out<=0;
   14284: out<=1;
   14285: out<=1;
   14286: out<=0;
   14287: out<=0;
   14288: out<=0;
   14289: out<=1;
   14290: out<=1;
   14291: out<=0;
   14292: out<=1;
   14293: out<=1;
   14294: out<=1;
   14295: out<=1;
   14296: out<=1;
   14297: out<=1;
   14298: out<=0;
   14299: out<=0;
   14300: out<=0;
   14301: out<=1;
   14302: out<=0;
   14303: out<=1;
   14304: out<=1;
   14305: out<=0;
   14306: out<=1;
   14307: out<=0;
   14308: out<=0;
   14309: out<=0;
   14310: out<=1;
   14311: out<=1;
   14312: out<=1;
   14313: out<=1;
   14314: out<=1;
   14315: out<=1;
   14316: out<=0;
   14317: out<=1;
   14318: out<=1;
   14319: out<=0;
   14320: out<=0;
   14321: out<=0;
   14322: out<=1;
   14323: out<=1;
   14324: out<=0;
   14325: out<=1;
   14326: out<=0;
   14327: out<=1;
   14328: out<=1;
   14329: out<=0;
   14330: out<=0;
   14331: out<=1;
   14332: out<=1;
   14333: out<=1;
   14334: out<=1;
   14335: out<=1;
   14336: out<=1;
   14337: out<=1;
   14338: out<=1;
   14339: out<=1;
   14340: out<=1;
   14341: out<=0;
   14342: out<=0;
   14343: out<=1;
   14344: out<=0;
   14345: out<=1;
   14346: out<=0;
   14347: out<=1;
   14348: out<=0;
   14349: out<=0;
   14350: out<=1;
   14351: out<=1;
   14352: out<=0;
   14353: out<=1;
   14354: out<=1;
   14355: out<=0;
   14356: out<=1;
   14357: out<=1;
   14358: out<=1;
   14359: out<=1;
   14360: out<=0;
   14361: out<=0;
   14362: out<=1;
   14363: out<=1;
   14364: out<=1;
   14365: out<=0;
   14366: out<=1;
   14367: out<=0;
   14368: out<=1;
   14369: out<=0;
   14370: out<=1;
   14371: out<=0;
   14372: out<=0;
   14373: out<=0;
   14374: out<=1;
   14375: out<=1;
   14376: out<=0;
   14377: out<=0;
   14378: out<=0;
   14379: out<=0;
   14380: out<=1;
   14381: out<=0;
   14382: out<=0;
   14383: out<=1;
   14384: out<=0;
   14385: out<=0;
   14386: out<=1;
   14387: out<=1;
   14388: out<=0;
   14389: out<=1;
   14390: out<=0;
   14391: out<=1;
   14392: out<=0;
   14393: out<=1;
   14394: out<=1;
   14395: out<=0;
   14396: out<=0;
   14397: out<=0;
   14398: out<=0;
   14399: out<=0;
   14400: out<=1;
   14401: out<=1;
   14402: out<=1;
   14403: out<=1;
   14404: out<=1;
   14405: out<=0;
   14406: out<=0;
   14407: out<=1;
   14408: out<=0;
   14409: out<=1;
   14410: out<=0;
   14411: out<=1;
   14412: out<=0;
   14413: out<=0;
   14414: out<=1;
   14415: out<=1;
   14416: out<=1;
   14417: out<=0;
   14418: out<=0;
   14419: out<=1;
   14420: out<=0;
   14421: out<=0;
   14422: out<=0;
   14423: out<=0;
   14424: out<=1;
   14425: out<=1;
   14426: out<=0;
   14427: out<=0;
   14428: out<=0;
   14429: out<=1;
   14430: out<=0;
   14431: out<=1;
   14432: out<=0;
   14433: out<=1;
   14434: out<=0;
   14435: out<=1;
   14436: out<=1;
   14437: out<=1;
   14438: out<=0;
   14439: out<=0;
   14440: out<=1;
   14441: out<=1;
   14442: out<=1;
   14443: out<=1;
   14444: out<=0;
   14445: out<=1;
   14446: out<=1;
   14447: out<=0;
   14448: out<=0;
   14449: out<=0;
   14450: out<=1;
   14451: out<=1;
   14452: out<=0;
   14453: out<=1;
   14454: out<=0;
   14455: out<=1;
   14456: out<=0;
   14457: out<=1;
   14458: out<=1;
   14459: out<=0;
   14460: out<=0;
   14461: out<=0;
   14462: out<=0;
   14463: out<=0;
   14464: out<=1;
   14465: out<=1;
   14466: out<=1;
   14467: out<=1;
   14468: out<=1;
   14469: out<=0;
   14470: out<=0;
   14471: out<=1;
   14472: out<=0;
   14473: out<=1;
   14474: out<=0;
   14475: out<=1;
   14476: out<=0;
   14477: out<=0;
   14478: out<=1;
   14479: out<=1;
   14480: out<=1;
   14481: out<=0;
   14482: out<=0;
   14483: out<=1;
   14484: out<=0;
   14485: out<=0;
   14486: out<=0;
   14487: out<=0;
   14488: out<=1;
   14489: out<=1;
   14490: out<=0;
   14491: out<=0;
   14492: out<=0;
   14493: out<=1;
   14494: out<=0;
   14495: out<=1;
   14496: out<=1;
   14497: out<=0;
   14498: out<=1;
   14499: out<=0;
   14500: out<=0;
   14501: out<=0;
   14502: out<=1;
   14503: out<=1;
   14504: out<=0;
   14505: out<=0;
   14506: out<=0;
   14507: out<=0;
   14508: out<=1;
   14509: out<=0;
   14510: out<=0;
   14511: out<=1;
   14512: out<=1;
   14513: out<=1;
   14514: out<=0;
   14515: out<=0;
   14516: out<=1;
   14517: out<=0;
   14518: out<=1;
   14519: out<=0;
   14520: out<=1;
   14521: out<=0;
   14522: out<=0;
   14523: out<=1;
   14524: out<=1;
   14525: out<=1;
   14526: out<=1;
   14527: out<=1;
   14528: out<=1;
   14529: out<=1;
   14530: out<=1;
   14531: out<=1;
   14532: out<=1;
   14533: out<=0;
   14534: out<=0;
   14535: out<=1;
   14536: out<=0;
   14537: out<=1;
   14538: out<=0;
   14539: out<=1;
   14540: out<=0;
   14541: out<=0;
   14542: out<=1;
   14543: out<=1;
   14544: out<=0;
   14545: out<=1;
   14546: out<=1;
   14547: out<=0;
   14548: out<=1;
   14549: out<=1;
   14550: out<=1;
   14551: out<=1;
   14552: out<=0;
   14553: out<=0;
   14554: out<=1;
   14555: out<=1;
   14556: out<=1;
   14557: out<=0;
   14558: out<=1;
   14559: out<=0;
   14560: out<=0;
   14561: out<=1;
   14562: out<=0;
   14563: out<=1;
   14564: out<=1;
   14565: out<=1;
   14566: out<=0;
   14567: out<=0;
   14568: out<=1;
   14569: out<=1;
   14570: out<=1;
   14571: out<=1;
   14572: out<=0;
   14573: out<=1;
   14574: out<=1;
   14575: out<=0;
   14576: out<=1;
   14577: out<=1;
   14578: out<=0;
   14579: out<=0;
   14580: out<=1;
   14581: out<=0;
   14582: out<=1;
   14583: out<=0;
   14584: out<=1;
   14585: out<=0;
   14586: out<=0;
   14587: out<=1;
   14588: out<=1;
   14589: out<=1;
   14590: out<=1;
   14591: out<=1;
   14592: out<=1;
   14593: out<=0;
   14594: out<=0;
   14595: out<=1;
   14596: out<=0;
   14597: out<=0;
   14598: out<=0;
   14599: out<=0;
   14600: out<=1;
   14601: out<=1;
   14602: out<=0;
   14603: out<=0;
   14604: out<=0;
   14605: out<=1;
   14606: out<=0;
   14607: out<=1;
   14608: out<=1;
   14609: out<=1;
   14610: out<=1;
   14611: out<=1;
   14612: out<=1;
   14613: out<=0;
   14614: out<=0;
   14615: out<=1;
   14616: out<=0;
   14617: out<=1;
   14618: out<=0;
   14619: out<=1;
   14620: out<=0;
   14621: out<=0;
   14622: out<=1;
   14623: out<=1;
   14624: out<=0;
   14625: out<=0;
   14626: out<=1;
   14627: out<=1;
   14628: out<=0;
   14629: out<=1;
   14630: out<=0;
   14631: out<=1;
   14632: out<=0;
   14633: out<=1;
   14634: out<=1;
   14635: out<=0;
   14636: out<=0;
   14637: out<=0;
   14638: out<=0;
   14639: out<=0;
   14640: out<=0;
   14641: out<=1;
   14642: out<=0;
   14643: out<=1;
   14644: out<=1;
   14645: out<=1;
   14646: out<=0;
   14647: out<=0;
   14648: out<=1;
   14649: out<=1;
   14650: out<=1;
   14651: out<=1;
   14652: out<=0;
   14653: out<=1;
   14654: out<=1;
   14655: out<=0;
   14656: out<=0;
   14657: out<=1;
   14658: out<=1;
   14659: out<=0;
   14660: out<=1;
   14661: out<=1;
   14662: out<=1;
   14663: out<=1;
   14664: out<=0;
   14665: out<=0;
   14666: out<=1;
   14667: out<=1;
   14668: out<=1;
   14669: out<=0;
   14670: out<=1;
   14671: out<=0;
   14672: out<=1;
   14673: out<=1;
   14674: out<=1;
   14675: out<=1;
   14676: out<=1;
   14677: out<=0;
   14678: out<=0;
   14679: out<=1;
   14680: out<=0;
   14681: out<=1;
   14682: out<=0;
   14683: out<=1;
   14684: out<=0;
   14685: out<=0;
   14686: out<=1;
   14687: out<=1;
   14688: out<=0;
   14689: out<=0;
   14690: out<=1;
   14691: out<=1;
   14692: out<=0;
   14693: out<=1;
   14694: out<=0;
   14695: out<=1;
   14696: out<=0;
   14697: out<=1;
   14698: out<=1;
   14699: out<=0;
   14700: out<=0;
   14701: out<=0;
   14702: out<=0;
   14703: out<=0;
   14704: out<=1;
   14705: out<=0;
   14706: out<=1;
   14707: out<=0;
   14708: out<=0;
   14709: out<=0;
   14710: out<=1;
   14711: out<=1;
   14712: out<=0;
   14713: out<=0;
   14714: out<=0;
   14715: out<=0;
   14716: out<=1;
   14717: out<=0;
   14718: out<=0;
   14719: out<=1;
   14720: out<=0;
   14721: out<=1;
   14722: out<=1;
   14723: out<=0;
   14724: out<=1;
   14725: out<=1;
   14726: out<=1;
   14727: out<=1;
   14728: out<=0;
   14729: out<=0;
   14730: out<=1;
   14731: out<=1;
   14732: out<=1;
   14733: out<=0;
   14734: out<=1;
   14735: out<=0;
   14736: out<=1;
   14737: out<=1;
   14738: out<=1;
   14739: out<=1;
   14740: out<=1;
   14741: out<=0;
   14742: out<=0;
   14743: out<=1;
   14744: out<=0;
   14745: out<=1;
   14746: out<=0;
   14747: out<=1;
   14748: out<=0;
   14749: out<=0;
   14750: out<=1;
   14751: out<=1;
   14752: out<=1;
   14753: out<=1;
   14754: out<=0;
   14755: out<=0;
   14756: out<=1;
   14757: out<=0;
   14758: out<=1;
   14759: out<=0;
   14760: out<=1;
   14761: out<=0;
   14762: out<=0;
   14763: out<=1;
   14764: out<=1;
   14765: out<=1;
   14766: out<=1;
   14767: out<=1;
   14768: out<=0;
   14769: out<=1;
   14770: out<=0;
   14771: out<=1;
   14772: out<=1;
   14773: out<=1;
   14774: out<=0;
   14775: out<=0;
   14776: out<=1;
   14777: out<=1;
   14778: out<=1;
   14779: out<=1;
   14780: out<=0;
   14781: out<=1;
   14782: out<=1;
   14783: out<=0;
   14784: out<=1;
   14785: out<=0;
   14786: out<=0;
   14787: out<=1;
   14788: out<=0;
   14789: out<=0;
   14790: out<=0;
   14791: out<=0;
   14792: out<=1;
   14793: out<=1;
   14794: out<=0;
   14795: out<=0;
   14796: out<=0;
   14797: out<=1;
   14798: out<=0;
   14799: out<=1;
   14800: out<=1;
   14801: out<=1;
   14802: out<=1;
   14803: out<=1;
   14804: out<=1;
   14805: out<=0;
   14806: out<=0;
   14807: out<=1;
   14808: out<=0;
   14809: out<=1;
   14810: out<=0;
   14811: out<=1;
   14812: out<=0;
   14813: out<=0;
   14814: out<=1;
   14815: out<=1;
   14816: out<=1;
   14817: out<=1;
   14818: out<=0;
   14819: out<=0;
   14820: out<=1;
   14821: out<=0;
   14822: out<=1;
   14823: out<=0;
   14824: out<=1;
   14825: out<=0;
   14826: out<=0;
   14827: out<=1;
   14828: out<=1;
   14829: out<=1;
   14830: out<=1;
   14831: out<=1;
   14832: out<=1;
   14833: out<=0;
   14834: out<=1;
   14835: out<=0;
   14836: out<=0;
   14837: out<=0;
   14838: out<=1;
   14839: out<=1;
   14840: out<=0;
   14841: out<=0;
   14842: out<=0;
   14843: out<=0;
   14844: out<=1;
   14845: out<=0;
   14846: out<=0;
   14847: out<=1;
   14848: out<=1;
   14849: out<=0;
   14850: out<=1;
   14851: out<=0;
   14852: out<=0;
   14853: out<=0;
   14854: out<=1;
   14855: out<=1;
   14856: out<=0;
   14857: out<=0;
   14858: out<=0;
   14859: out<=0;
   14860: out<=1;
   14861: out<=0;
   14862: out<=0;
   14863: out<=1;
   14864: out<=1;
   14865: out<=1;
   14866: out<=0;
   14867: out<=0;
   14868: out<=1;
   14869: out<=0;
   14870: out<=1;
   14871: out<=0;
   14872: out<=1;
   14873: out<=0;
   14874: out<=0;
   14875: out<=1;
   14876: out<=1;
   14877: out<=1;
   14878: out<=1;
   14879: out<=1;
   14880: out<=1;
   14881: out<=1;
   14882: out<=1;
   14883: out<=1;
   14884: out<=1;
   14885: out<=0;
   14886: out<=0;
   14887: out<=1;
   14888: out<=0;
   14889: out<=1;
   14890: out<=0;
   14891: out<=1;
   14892: out<=0;
   14893: out<=0;
   14894: out<=1;
   14895: out<=1;
   14896: out<=1;
   14897: out<=0;
   14898: out<=0;
   14899: out<=1;
   14900: out<=0;
   14901: out<=0;
   14902: out<=0;
   14903: out<=0;
   14904: out<=1;
   14905: out<=1;
   14906: out<=0;
   14907: out<=0;
   14908: out<=0;
   14909: out<=1;
   14910: out<=0;
   14911: out<=1;
   14912: out<=0;
   14913: out<=1;
   14914: out<=0;
   14915: out<=1;
   14916: out<=1;
   14917: out<=1;
   14918: out<=0;
   14919: out<=0;
   14920: out<=1;
   14921: out<=1;
   14922: out<=1;
   14923: out<=1;
   14924: out<=0;
   14925: out<=1;
   14926: out<=1;
   14927: out<=0;
   14928: out<=1;
   14929: out<=1;
   14930: out<=0;
   14931: out<=0;
   14932: out<=1;
   14933: out<=0;
   14934: out<=1;
   14935: out<=0;
   14936: out<=1;
   14937: out<=0;
   14938: out<=0;
   14939: out<=1;
   14940: out<=1;
   14941: out<=1;
   14942: out<=1;
   14943: out<=1;
   14944: out<=1;
   14945: out<=1;
   14946: out<=1;
   14947: out<=1;
   14948: out<=1;
   14949: out<=0;
   14950: out<=0;
   14951: out<=1;
   14952: out<=0;
   14953: out<=1;
   14954: out<=0;
   14955: out<=1;
   14956: out<=0;
   14957: out<=0;
   14958: out<=1;
   14959: out<=1;
   14960: out<=0;
   14961: out<=1;
   14962: out<=1;
   14963: out<=0;
   14964: out<=1;
   14965: out<=1;
   14966: out<=1;
   14967: out<=1;
   14968: out<=0;
   14969: out<=0;
   14970: out<=1;
   14971: out<=1;
   14972: out<=1;
   14973: out<=0;
   14974: out<=1;
   14975: out<=0;
   14976: out<=1;
   14977: out<=0;
   14978: out<=1;
   14979: out<=0;
   14980: out<=0;
   14981: out<=0;
   14982: out<=1;
   14983: out<=1;
   14984: out<=0;
   14985: out<=0;
   14986: out<=0;
   14987: out<=0;
   14988: out<=1;
   14989: out<=0;
   14990: out<=0;
   14991: out<=1;
   14992: out<=0;
   14993: out<=0;
   14994: out<=1;
   14995: out<=1;
   14996: out<=0;
   14997: out<=1;
   14998: out<=0;
   14999: out<=1;
   15000: out<=0;
   15001: out<=1;
   15002: out<=1;
   15003: out<=0;
   15004: out<=0;
   15005: out<=0;
   15006: out<=0;
   15007: out<=0;
   15008: out<=1;
   15009: out<=1;
   15010: out<=1;
   15011: out<=1;
   15012: out<=1;
   15013: out<=0;
   15014: out<=0;
   15015: out<=1;
   15016: out<=0;
   15017: out<=1;
   15018: out<=0;
   15019: out<=1;
   15020: out<=0;
   15021: out<=0;
   15022: out<=1;
   15023: out<=1;
   15024: out<=0;
   15025: out<=1;
   15026: out<=1;
   15027: out<=0;
   15028: out<=1;
   15029: out<=1;
   15030: out<=1;
   15031: out<=1;
   15032: out<=0;
   15033: out<=0;
   15034: out<=1;
   15035: out<=1;
   15036: out<=1;
   15037: out<=0;
   15038: out<=1;
   15039: out<=0;
   15040: out<=0;
   15041: out<=1;
   15042: out<=0;
   15043: out<=1;
   15044: out<=1;
   15045: out<=1;
   15046: out<=0;
   15047: out<=0;
   15048: out<=1;
   15049: out<=1;
   15050: out<=1;
   15051: out<=1;
   15052: out<=0;
   15053: out<=1;
   15054: out<=1;
   15055: out<=0;
   15056: out<=0;
   15057: out<=0;
   15058: out<=1;
   15059: out<=1;
   15060: out<=0;
   15061: out<=1;
   15062: out<=0;
   15063: out<=1;
   15064: out<=0;
   15065: out<=1;
   15066: out<=1;
   15067: out<=0;
   15068: out<=0;
   15069: out<=0;
   15070: out<=0;
   15071: out<=0;
   15072: out<=1;
   15073: out<=1;
   15074: out<=1;
   15075: out<=1;
   15076: out<=1;
   15077: out<=0;
   15078: out<=0;
   15079: out<=1;
   15080: out<=0;
   15081: out<=1;
   15082: out<=0;
   15083: out<=1;
   15084: out<=0;
   15085: out<=0;
   15086: out<=1;
   15087: out<=1;
   15088: out<=1;
   15089: out<=0;
   15090: out<=0;
   15091: out<=1;
   15092: out<=0;
   15093: out<=0;
   15094: out<=0;
   15095: out<=0;
   15096: out<=1;
   15097: out<=1;
   15098: out<=0;
   15099: out<=0;
   15100: out<=0;
   15101: out<=1;
   15102: out<=0;
   15103: out<=1;
   15104: out<=1;
   15105: out<=1;
   15106: out<=0;
   15107: out<=0;
   15108: out<=1;
   15109: out<=0;
   15110: out<=1;
   15111: out<=0;
   15112: out<=1;
   15113: out<=0;
   15114: out<=0;
   15115: out<=1;
   15116: out<=1;
   15117: out<=1;
   15118: out<=1;
   15119: out<=1;
   15120: out<=0;
   15121: out<=1;
   15122: out<=0;
   15123: out<=1;
   15124: out<=1;
   15125: out<=1;
   15126: out<=0;
   15127: out<=0;
   15128: out<=1;
   15129: out<=1;
   15130: out<=1;
   15131: out<=1;
   15132: out<=0;
   15133: out<=1;
   15134: out<=1;
   15135: out<=0;
   15136: out<=0;
   15137: out<=1;
   15138: out<=1;
   15139: out<=0;
   15140: out<=1;
   15141: out<=1;
   15142: out<=1;
   15143: out<=1;
   15144: out<=0;
   15145: out<=0;
   15146: out<=1;
   15147: out<=1;
   15148: out<=1;
   15149: out<=0;
   15150: out<=1;
   15151: out<=0;
   15152: out<=1;
   15153: out<=1;
   15154: out<=1;
   15155: out<=1;
   15156: out<=1;
   15157: out<=0;
   15158: out<=0;
   15159: out<=1;
   15160: out<=0;
   15161: out<=1;
   15162: out<=0;
   15163: out<=1;
   15164: out<=0;
   15165: out<=0;
   15166: out<=1;
   15167: out<=1;
   15168: out<=1;
   15169: out<=1;
   15170: out<=0;
   15171: out<=0;
   15172: out<=1;
   15173: out<=0;
   15174: out<=1;
   15175: out<=0;
   15176: out<=1;
   15177: out<=0;
   15178: out<=0;
   15179: out<=1;
   15180: out<=1;
   15181: out<=1;
   15182: out<=1;
   15183: out<=1;
   15184: out<=1;
   15185: out<=0;
   15186: out<=1;
   15187: out<=0;
   15188: out<=0;
   15189: out<=0;
   15190: out<=1;
   15191: out<=1;
   15192: out<=0;
   15193: out<=0;
   15194: out<=0;
   15195: out<=0;
   15196: out<=1;
   15197: out<=0;
   15198: out<=0;
   15199: out<=1;
   15200: out<=1;
   15201: out<=0;
   15202: out<=0;
   15203: out<=1;
   15204: out<=0;
   15205: out<=0;
   15206: out<=0;
   15207: out<=0;
   15208: out<=1;
   15209: out<=1;
   15210: out<=0;
   15211: out<=0;
   15212: out<=0;
   15213: out<=1;
   15214: out<=0;
   15215: out<=1;
   15216: out<=1;
   15217: out<=1;
   15218: out<=1;
   15219: out<=1;
   15220: out<=1;
   15221: out<=0;
   15222: out<=0;
   15223: out<=1;
   15224: out<=0;
   15225: out<=1;
   15226: out<=0;
   15227: out<=1;
   15228: out<=0;
   15229: out<=0;
   15230: out<=1;
   15231: out<=1;
   15232: out<=0;
   15233: out<=0;
   15234: out<=1;
   15235: out<=1;
   15236: out<=0;
   15237: out<=1;
   15238: out<=0;
   15239: out<=1;
   15240: out<=0;
   15241: out<=1;
   15242: out<=1;
   15243: out<=0;
   15244: out<=0;
   15245: out<=0;
   15246: out<=0;
   15247: out<=0;
   15248: out<=0;
   15249: out<=1;
   15250: out<=0;
   15251: out<=1;
   15252: out<=1;
   15253: out<=1;
   15254: out<=0;
   15255: out<=0;
   15256: out<=1;
   15257: out<=1;
   15258: out<=1;
   15259: out<=1;
   15260: out<=0;
   15261: out<=1;
   15262: out<=1;
   15263: out<=0;
   15264: out<=1;
   15265: out<=0;
   15266: out<=0;
   15267: out<=1;
   15268: out<=0;
   15269: out<=0;
   15270: out<=0;
   15271: out<=0;
   15272: out<=1;
   15273: out<=1;
   15274: out<=0;
   15275: out<=0;
   15276: out<=0;
   15277: out<=1;
   15278: out<=0;
   15279: out<=1;
   15280: out<=1;
   15281: out<=1;
   15282: out<=1;
   15283: out<=1;
   15284: out<=1;
   15285: out<=0;
   15286: out<=0;
   15287: out<=1;
   15288: out<=0;
   15289: out<=1;
   15290: out<=0;
   15291: out<=1;
   15292: out<=0;
   15293: out<=0;
   15294: out<=1;
   15295: out<=1;
   15296: out<=0;
   15297: out<=0;
   15298: out<=1;
   15299: out<=1;
   15300: out<=0;
   15301: out<=1;
   15302: out<=0;
   15303: out<=1;
   15304: out<=0;
   15305: out<=1;
   15306: out<=1;
   15307: out<=0;
   15308: out<=0;
   15309: out<=0;
   15310: out<=0;
   15311: out<=0;
   15312: out<=1;
   15313: out<=0;
   15314: out<=1;
   15315: out<=0;
   15316: out<=0;
   15317: out<=0;
   15318: out<=1;
   15319: out<=1;
   15320: out<=0;
   15321: out<=0;
   15322: out<=0;
   15323: out<=0;
   15324: out<=1;
   15325: out<=0;
   15326: out<=0;
   15327: out<=1;
   15328: out<=0;
   15329: out<=1;
   15330: out<=1;
   15331: out<=0;
   15332: out<=1;
   15333: out<=1;
   15334: out<=1;
   15335: out<=1;
   15336: out<=0;
   15337: out<=0;
   15338: out<=1;
   15339: out<=1;
   15340: out<=1;
   15341: out<=0;
   15342: out<=1;
   15343: out<=0;
   15344: out<=1;
   15345: out<=1;
   15346: out<=1;
   15347: out<=1;
   15348: out<=1;
   15349: out<=0;
   15350: out<=0;
   15351: out<=1;
   15352: out<=0;
   15353: out<=1;
   15354: out<=0;
   15355: out<=1;
   15356: out<=0;
   15357: out<=0;
   15358: out<=1;
   15359: out<=1;
   15360: out<=0;
   15361: out<=1;
   15362: out<=1;
   15363: out<=0;
   15364: out<=0;
   15365: out<=0;
   15366: out<=0;
   15367: out<=0;
   15368: out<=1;
   15369: out<=1;
   15370: out<=0;
   15371: out<=0;
   15372: out<=1;
   15373: out<=0;
   15374: out<=1;
   15375: out<=0;
   15376: out<=1;
   15377: out<=1;
   15378: out<=1;
   15379: out<=1;
   15380: out<=0;
   15381: out<=1;
   15382: out<=1;
   15383: out<=0;
   15384: out<=1;
   15385: out<=0;
   15386: out<=1;
   15387: out<=0;
   15388: out<=0;
   15389: out<=0;
   15390: out<=1;
   15391: out<=1;
   15392: out<=0;
   15393: out<=0;
   15394: out<=1;
   15395: out<=1;
   15396: out<=1;
   15397: out<=0;
   15398: out<=1;
   15399: out<=0;
   15400: out<=1;
   15401: out<=0;
   15402: out<=0;
   15403: out<=1;
   15404: out<=0;
   15405: out<=0;
   15406: out<=0;
   15407: out<=0;
   15408: out<=1;
   15409: out<=0;
   15410: out<=1;
   15411: out<=0;
   15412: out<=1;
   15413: out<=1;
   15414: out<=0;
   15415: out<=0;
   15416: out<=1;
   15417: out<=1;
   15418: out<=1;
   15419: out<=1;
   15420: out<=1;
   15421: out<=0;
   15422: out<=0;
   15423: out<=1;
   15424: out<=1;
   15425: out<=0;
   15426: out<=0;
   15427: out<=1;
   15428: out<=1;
   15429: out<=1;
   15430: out<=1;
   15431: out<=1;
   15432: out<=0;
   15433: out<=0;
   15434: out<=1;
   15435: out<=1;
   15436: out<=0;
   15437: out<=1;
   15438: out<=0;
   15439: out<=1;
   15440: out<=1;
   15441: out<=1;
   15442: out<=1;
   15443: out<=1;
   15444: out<=0;
   15445: out<=1;
   15446: out<=1;
   15447: out<=0;
   15448: out<=1;
   15449: out<=0;
   15450: out<=1;
   15451: out<=0;
   15452: out<=0;
   15453: out<=0;
   15454: out<=1;
   15455: out<=1;
   15456: out<=0;
   15457: out<=0;
   15458: out<=1;
   15459: out<=1;
   15460: out<=1;
   15461: out<=0;
   15462: out<=1;
   15463: out<=0;
   15464: out<=1;
   15465: out<=0;
   15466: out<=0;
   15467: out<=1;
   15468: out<=0;
   15469: out<=0;
   15470: out<=0;
   15471: out<=0;
   15472: out<=0;
   15473: out<=1;
   15474: out<=0;
   15475: out<=1;
   15476: out<=0;
   15477: out<=0;
   15478: out<=1;
   15479: out<=1;
   15480: out<=0;
   15481: out<=0;
   15482: out<=0;
   15483: out<=0;
   15484: out<=0;
   15485: out<=1;
   15486: out<=1;
   15487: out<=0;
   15488: out<=1;
   15489: out<=0;
   15490: out<=0;
   15491: out<=1;
   15492: out<=1;
   15493: out<=1;
   15494: out<=1;
   15495: out<=1;
   15496: out<=0;
   15497: out<=0;
   15498: out<=1;
   15499: out<=1;
   15500: out<=0;
   15501: out<=1;
   15502: out<=0;
   15503: out<=1;
   15504: out<=1;
   15505: out<=1;
   15506: out<=1;
   15507: out<=1;
   15508: out<=0;
   15509: out<=1;
   15510: out<=1;
   15511: out<=0;
   15512: out<=1;
   15513: out<=0;
   15514: out<=1;
   15515: out<=0;
   15516: out<=0;
   15517: out<=0;
   15518: out<=1;
   15519: out<=1;
   15520: out<=1;
   15521: out<=1;
   15522: out<=0;
   15523: out<=0;
   15524: out<=0;
   15525: out<=1;
   15526: out<=0;
   15527: out<=1;
   15528: out<=0;
   15529: out<=1;
   15530: out<=1;
   15531: out<=0;
   15532: out<=1;
   15533: out<=1;
   15534: out<=1;
   15535: out<=1;
   15536: out<=1;
   15537: out<=0;
   15538: out<=1;
   15539: out<=0;
   15540: out<=1;
   15541: out<=1;
   15542: out<=0;
   15543: out<=0;
   15544: out<=1;
   15545: out<=1;
   15546: out<=1;
   15547: out<=1;
   15548: out<=1;
   15549: out<=0;
   15550: out<=0;
   15551: out<=1;
   15552: out<=0;
   15553: out<=1;
   15554: out<=1;
   15555: out<=0;
   15556: out<=0;
   15557: out<=0;
   15558: out<=0;
   15559: out<=0;
   15560: out<=1;
   15561: out<=1;
   15562: out<=0;
   15563: out<=0;
   15564: out<=1;
   15565: out<=0;
   15566: out<=1;
   15567: out<=0;
   15568: out<=1;
   15569: out<=1;
   15570: out<=1;
   15571: out<=1;
   15572: out<=0;
   15573: out<=1;
   15574: out<=1;
   15575: out<=0;
   15576: out<=1;
   15577: out<=0;
   15578: out<=1;
   15579: out<=0;
   15580: out<=0;
   15581: out<=0;
   15582: out<=1;
   15583: out<=1;
   15584: out<=1;
   15585: out<=1;
   15586: out<=0;
   15587: out<=0;
   15588: out<=0;
   15589: out<=1;
   15590: out<=0;
   15591: out<=1;
   15592: out<=0;
   15593: out<=1;
   15594: out<=1;
   15595: out<=0;
   15596: out<=1;
   15597: out<=1;
   15598: out<=1;
   15599: out<=1;
   15600: out<=0;
   15601: out<=1;
   15602: out<=0;
   15603: out<=1;
   15604: out<=0;
   15605: out<=0;
   15606: out<=1;
   15607: out<=1;
   15608: out<=0;
   15609: out<=0;
   15610: out<=0;
   15611: out<=0;
   15612: out<=0;
   15613: out<=1;
   15614: out<=1;
   15615: out<=0;
   15616: out<=1;
   15617: out<=1;
   15618: out<=1;
   15619: out<=1;
   15620: out<=0;
   15621: out<=1;
   15622: out<=1;
   15623: out<=0;
   15624: out<=1;
   15625: out<=0;
   15626: out<=1;
   15627: out<=0;
   15628: out<=0;
   15629: out<=0;
   15630: out<=1;
   15631: out<=1;
   15632: out<=1;
   15633: out<=0;
   15634: out<=0;
   15635: out<=1;
   15636: out<=1;
   15637: out<=1;
   15638: out<=1;
   15639: out<=1;
   15640: out<=0;
   15641: out<=0;
   15642: out<=1;
   15643: out<=1;
   15644: out<=0;
   15645: out<=1;
   15646: out<=0;
   15647: out<=1;
   15648: out<=0;
   15649: out<=1;
   15650: out<=0;
   15651: out<=1;
   15652: out<=0;
   15653: out<=0;
   15654: out<=1;
   15655: out<=1;
   15656: out<=0;
   15657: out<=0;
   15658: out<=0;
   15659: out<=0;
   15660: out<=0;
   15661: out<=1;
   15662: out<=1;
   15663: out<=0;
   15664: out<=0;
   15665: out<=0;
   15666: out<=1;
   15667: out<=1;
   15668: out<=1;
   15669: out<=0;
   15670: out<=1;
   15671: out<=0;
   15672: out<=1;
   15673: out<=0;
   15674: out<=0;
   15675: out<=1;
   15676: out<=0;
   15677: out<=0;
   15678: out<=0;
   15679: out<=0;
   15680: out<=1;
   15681: out<=1;
   15682: out<=1;
   15683: out<=1;
   15684: out<=0;
   15685: out<=1;
   15686: out<=1;
   15687: out<=0;
   15688: out<=1;
   15689: out<=0;
   15690: out<=1;
   15691: out<=0;
   15692: out<=0;
   15693: out<=0;
   15694: out<=1;
   15695: out<=1;
   15696: out<=0;
   15697: out<=1;
   15698: out<=1;
   15699: out<=0;
   15700: out<=0;
   15701: out<=0;
   15702: out<=0;
   15703: out<=0;
   15704: out<=1;
   15705: out<=1;
   15706: out<=0;
   15707: out<=0;
   15708: out<=1;
   15709: out<=0;
   15710: out<=1;
   15711: out<=0;
   15712: out<=1;
   15713: out<=0;
   15714: out<=1;
   15715: out<=0;
   15716: out<=1;
   15717: out<=1;
   15718: out<=0;
   15719: out<=0;
   15720: out<=1;
   15721: out<=1;
   15722: out<=1;
   15723: out<=1;
   15724: out<=1;
   15725: out<=0;
   15726: out<=0;
   15727: out<=1;
   15728: out<=0;
   15729: out<=0;
   15730: out<=1;
   15731: out<=1;
   15732: out<=1;
   15733: out<=0;
   15734: out<=1;
   15735: out<=0;
   15736: out<=1;
   15737: out<=0;
   15738: out<=0;
   15739: out<=1;
   15740: out<=0;
   15741: out<=0;
   15742: out<=0;
   15743: out<=0;
   15744: out<=1;
   15745: out<=1;
   15746: out<=1;
   15747: out<=1;
   15748: out<=0;
   15749: out<=1;
   15750: out<=1;
   15751: out<=0;
   15752: out<=1;
   15753: out<=0;
   15754: out<=1;
   15755: out<=0;
   15756: out<=0;
   15757: out<=0;
   15758: out<=1;
   15759: out<=1;
   15760: out<=0;
   15761: out<=1;
   15762: out<=1;
   15763: out<=0;
   15764: out<=0;
   15765: out<=0;
   15766: out<=0;
   15767: out<=0;
   15768: out<=1;
   15769: out<=1;
   15770: out<=0;
   15771: out<=0;
   15772: out<=1;
   15773: out<=0;
   15774: out<=1;
   15775: out<=0;
   15776: out<=0;
   15777: out<=1;
   15778: out<=0;
   15779: out<=1;
   15780: out<=0;
   15781: out<=0;
   15782: out<=1;
   15783: out<=1;
   15784: out<=0;
   15785: out<=0;
   15786: out<=0;
   15787: out<=0;
   15788: out<=0;
   15789: out<=1;
   15790: out<=1;
   15791: out<=0;
   15792: out<=1;
   15793: out<=1;
   15794: out<=0;
   15795: out<=0;
   15796: out<=0;
   15797: out<=1;
   15798: out<=0;
   15799: out<=1;
   15800: out<=0;
   15801: out<=1;
   15802: out<=1;
   15803: out<=0;
   15804: out<=1;
   15805: out<=1;
   15806: out<=1;
   15807: out<=1;
   15808: out<=1;
   15809: out<=1;
   15810: out<=1;
   15811: out<=1;
   15812: out<=0;
   15813: out<=1;
   15814: out<=1;
   15815: out<=0;
   15816: out<=1;
   15817: out<=0;
   15818: out<=1;
   15819: out<=0;
   15820: out<=0;
   15821: out<=0;
   15822: out<=1;
   15823: out<=1;
   15824: out<=1;
   15825: out<=0;
   15826: out<=0;
   15827: out<=1;
   15828: out<=1;
   15829: out<=1;
   15830: out<=1;
   15831: out<=1;
   15832: out<=0;
   15833: out<=0;
   15834: out<=1;
   15835: out<=1;
   15836: out<=0;
   15837: out<=1;
   15838: out<=0;
   15839: out<=1;
   15840: out<=1;
   15841: out<=0;
   15842: out<=1;
   15843: out<=0;
   15844: out<=1;
   15845: out<=1;
   15846: out<=0;
   15847: out<=0;
   15848: out<=1;
   15849: out<=1;
   15850: out<=1;
   15851: out<=1;
   15852: out<=1;
   15853: out<=0;
   15854: out<=0;
   15855: out<=1;
   15856: out<=1;
   15857: out<=1;
   15858: out<=0;
   15859: out<=0;
   15860: out<=0;
   15861: out<=1;
   15862: out<=0;
   15863: out<=1;
   15864: out<=0;
   15865: out<=1;
   15866: out<=1;
   15867: out<=0;
   15868: out<=1;
   15869: out<=1;
   15870: out<=1;
   15871: out<=1;
   15872: out<=1;
   15873: out<=1;
   15874: out<=0;
   15875: out<=0;
   15876: out<=0;
   15877: out<=1;
   15878: out<=0;
   15879: out<=1;
   15880: out<=0;
   15881: out<=1;
   15882: out<=1;
   15883: out<=0;
   15884: out<=1;
   15885: out<=1;
   15886: out<=1;
   15887: out<=1;
   15888: out<=1;
   15889: out<=0;
   15890: out<=1;
   15891: out<=0;
   15892: out<=1;
   15893: out<=1;
   15894: out<=0;
   15895: out<=0;
   15896: out<=1;
   15897: out<=1;
   15898: out<=1;
   15899: out<=1;
   15900: out<=1;
   15901: out<=0;
   15902: out<=0;
   15903: out<=1;
   15904: out<=1;
   15905: out<=0;
   15906: out<=0;
   15907: out<=1;
   15908: out<=1;
   15909: out<=1;
   15910: out<=1;
   15911: out<=1;
   15912: out<=0;
   15913: out<=0;
   15914: out<=1;
   15915: out<=1;
   15916: out<=0;
   15917: out<=1;
   15918: out<=0;
   15919: out<=1;
   15920: out<=1;
   15921: out<=1;
   15922: out<=1;
   15923: out<=1;
   15924: out<=0;
   15925: out<=1;
   15926: out<=1;
   15927: out<=0;
   15928: out<=1;
   15929: out<=0;
   15930: out<=1;
   15931: out<=0;
   15932: out<=0;
   15933: out<=0;
   15934: out<=1;
   15935: out<=1;
   15936: out<=1;
   15937: out<=1;
   15938: out<=0;
   15939: out<=0;
   15940: out<=0;
   15941: out<=1;
   15942: out<=0;
   15943: out<=1;
   15944: out<=0;
   15945: out<=1;
   15946: out<=1;
   15947: out<=0;
   15948: out<=1;
   15949: out<=1;
   15950: out<=1;
   15951: out<=1;
   15952: out<=0;
   15953: out<=1;
   15954: out<=0;
   15955: out<=1;
   15956: out<=0;
   15957: out<=0;
   15958: out<=1;
   15959: out<=1;
   15960: out<=0;
   15961: out<=0;
   15962: out<=0;
   15963: out<=0;
   15964: out<=0;
   15965: out<=1;
   15966: out<=1;
   15967: out<=0;
   15968: out<=0;
   15969: out<=1;
   15970: out<=1;
   15971: out<=0;
   15972: out<=0;
   15973: out<=0;
   15974: out<=0;
   15975: out<=0;
   15976: out<=1;
   15977: out<=1;
   15978: out<=0;
   15979: out<=0;
   15980: out<=1;
   15981: out<=0;
   15982: out<=1;
   15983: out<=0;
   15984: out<=1;
   15985: out<=1;
   15986: out<=1;
   15987: out<=1;
   15988: out<=0;
   15989: out<=1;
   15990: out<=1;
   15991: out<=0;
   15992: out<=1;
   15993: out<=0;
   15994: out<=1;
   15995: out<=0;
   15996: out<=0;
   15997: out<=0;
   15998: out<=1;
   15999: out<=1;
   16000: out<=0;
   16001: out<=0;
   16002: out<=1;
   16003: out<=1;
   16004: out<=1;
   16005: out<=0;
   16006: out<=1;
   16007: out<=0;
   16008: out<=1;
   16009: out<=0;
   16010: out<=0;
   16011: out<=1;
   16012: out<=0;
   16013: out<=0;
   16014: out<=0;
   16015: out<=0;
   16016: out<=1;
   16017: out<=0;
   16018: out<=1;
   16019: out<=0;
   16020: out<=1;
   16021: out<=1;
   16022: out<=0;
   16023: out<=0;
   16024: out<=1;
   16025: out<=1;
   16026: out<=1;
   16027: out<=1;
   16028: out<=1;
   16029: out<=0;
   16030: out<=0;
   16031: out<=1;
   16032: out<=0;
   16033: out<=1;
   16034: out<=1;
   16035: out<=0;
   16036: out<=0;
   16037: out<=0;
   16038: out<=0;
   16039: out<=0;
   16040: out<=1;
   16041: out<=1;
   16042: out<=0;
   16043: out<=0;
   16044: out<=1;
   16045: out<=0;
   16046: out<=1;
   16047: out<=0;
   16048: out<=1;
   16049: out<=1;
   16050: out<=1;
   16051: out<=1;
   16052: out<=0;
   16053: out<=1;
   16054: out<=1;
   16055: out<=0;
   16056: out<=1;
   16057: out<=0;
   16058: out<=1;
   16059: out<=0;
   16060: out<=0;
   16061: out<=0;
   16062: out<=1;
   16063: out<=1;
   16064: out<=0;
   16065: out<=0;
   16066: out<=1;
   16067: out<=1;
   16068: out<=1;
   16069: out<=0;
   16070: out<=1;
   16071: out<=0;
   16072: out<=1;
   16073: out<=0;
   16074: out<=0;
   16075: out<=1;
   16076: out<=0;
   16077: out<=0;
   16078: out<=0;
   16079: out<=0;
   16080: out<=0;
   16081: out<=1;
   16082: out<=0;
   16083: out<=1;
   16084: out<=0;
   16085: out<=0;
   16086: out<=1;
   16087: out<=1;
   16088: out<=0;
   16089: out<=0;
   16090: out<=0;
   16091: out<=0;
   16092: out<=0;
   16093: out<=1;
   16094: out<=1;
   16095: out<=0;
   16096: out<=1;
   16097: out<=0;
   16098: out<=0;
   16099: out<=1;
   16100: out<=1;
   16101: out<=1;
   16102: out<=1;
   16103: out<=1;
   16104: out<=0;
   16105: out<=0;
   16106: out<=1;
   16107: out<=1;
   16108: out<=0;
   16109: out<=1;
   16110: out<=0;
   16111: out<=1;
   16112: out<=1;
   16113: out<=1;
   16114: out<=1;
   16115: out<=1;
   16116: out<=0;
   16117: out<=1;
   16118: out<=1;
   16119: out<=0;
   16120: out<=1;
   16121: out<=0;
   16122: out<=1;
   16123: out<=0;
   16124: out<=0;
   16125: out<=0;
   16126: out<=1;
   16127: out<=1;
   16128: out<=0;
   16129: out<=1;
   16130: out<=0;
   16131: out<=1;
   16132: out<=0;
   16133: out<=0;
   16134: out<=1;
   16135: out<=1;
   16136: out<=0;
   16137: out<=0;
   16138: out<=0;
   16139: out<=0;
   16140: out<=0;
   16141: out<=1;
   16142: out<=1;
   16143: out<=0;
   16144: out<=1;
   16145: out<=1;
   16146: out<=0;
   16147: out<=0;
   16148: out<=0;
   16149: out<=1;
   16150: out<=0;
   16151: out<=1;
   16152: out<=0;
   16153: out<=1;
   16154: out<=1;
   16155: out<=0;
   16156: out<=1;
   16157: out<=1;
   16158: out<=1;
   16159: out<=1;
   16160: out<=1;
   16161: out<=1;
   16162: out<=1;
   16163: out<=1;
   16164: out<=0;
   16165: out<=1;
   16166: out<=1;
   16167: out<=0;
   16168: out<=1;
   16169: out<=0;
   16170: out<=1;
   16171: out<=0;
   16172: out<=0;
   16173: out<=0;
   16174: out<=1;
   16175: out<=1;
   16176: out<=0;
   16177: out<=1;
   16178: out<=1;
   16179: out<=0;
   16180: out<=0;
   16181: out<=0;
   16182: out<=0;
   16183: out<=0;
   16184: out<=1;
   16185: out<=1;
   16186: out<=0;
   16187: out<=0;
   16188: out<=1;
   16189: out<=0;
   16190: out<=1;
   16191: out<=0;
   16192: out<=1;
   16193: out<=0;
   16194: out<=1;
   16195: out<=0;
   16196: out<=1;
   16197: out<=1;
   16198: out<=0;
   16199: out<=0;
   16200: out<=1;
   16201: out<=1;
   16202: out<=1;
   16203: out<=1;
   16204: out<=1;
   16205: out<=0;
   16206: out<=0;
   16207: out<=1;
   16208: out<=1;
   16209: out<=1;
   16210: out<=0;
   16211: out<=0;
   16212: out<=0;
   16213: out<=1;
   16214: out<=0;
   16215: out<=1;
   16216: out<=0;
   16217: out<=1;
   16218: out<=1;
   16219: out<=0;
   16220: out<=1;
   16221: out<=1;
   16222: out<=1;
   16223: out<=1;
   16224: out<=1;
   16225: out<=1;
   16226: out<=1;
   16227: out<=1;
   16228: out<=0;
   16229: out<=1;
   16230: out<=1;
   16231: out<=0;
   16232: out<=1;
   16233: out<=0;
   16234: out<=1;
   16235: out<=0;
   16236: out<=0;
   16237: out<=0;
   16238: out<=1;
   16239: out<=1;
   16240: out<=1;
   16241: out<=0;
   16242: out<=0;
   16243: out<=1;
   16244: out<=1;
   16245: out<=1;
   16246: out<=1;
   16247: out<=1;
   16248: out<=0;
   16249: out<=0;
   16250: out<=1;
   16251: out<=1;
   16252: out<=0;
   16253: out<=1;
   16254: out<=0;
   16255: out<=1;
   16256: out<=0;
   16257: out<=1;
   16258: out<=0;
   16259: out<=1;
   16260: out<=0;
   16261: out<=0;
   16262: out<=1;
   16263: out<=1;
   16264: out<=0;
   16265: out<=0;
   16266: out<=0;
   16267: out<=0;
   16268: out<=0;
   16269: out<=1;
   16270: out<=1;
   16271: out<=0;
   16272: out<=0;
   16273: out<=0;
   16274: out<=1;
   16275: out<=1;
   16276: out<=1;
   16277: out<=0;
   16278: out<=1;
   16279: out<=0;
   16280: out<=1;
   16281: out<=0;
   16282: out<=0;
   16283: out<=1;
   16284: out<=0;
   16285: out<=0;
   16286: out<=0;
   16287: out<=0;
   16288: out<=1;
   16289: out<=1;
   16290: out<=1;
   16291: out<=1;
   16292: out<=0;
   16293: out<=1;
   16294: out<=1;
   16295: out<=0;
   16296: out<=1;
   16297: out<=0;
   16298: out<=1;
   16299: out<=0;
   16300: out<=0;
   16301: out<=0;
   16302: out<=1;
   16303: out<=1;
   16304: out<=1;
   16305: out<=0;
   16306: out<=0;
   16307: out<=1;
   16308: out<=1;
   16309: out<=1;
   16310: out<=1;
   16311: out<=1;
   16312: out<=0;
   16313: out<=0;
   16314: out<=1;
   16315: out<=1;
   16316: out<=0;
   16317: out<=1;
   16318: out<=0;
   16319: out<=1;
   16320: out<=1;
   16321: out<=0;
   16322: out<=1;
   16323: out<=0;
   16324: out<=1;
   16325: out<=1;
   16326: out<=0;
   16327: out<=0;
   16328: out<=1;
   16329: out<=1;
   16330: out<=1;
   16331: out<=1;
   16332: out<=1;
   16333: out<=0;
   16334: out<=0;
   16335: out<=1;
   16336: out<=0;
   16337: out<=0;
   16338: out<=1;
   16339: out<=1;
   16340: out<=1;
   16341: out<=0;
   16342: out<=1;
   16343: out<=0;
   16344: out<=1;
   16345: out<=0;
   16346: out<=0;
   16347: out<=1;
   16348: out<=0;
   16349: out<=0;
   16350: out<=0;
   16351: out<=0;
   16352: out<=1;
   16353: out<=1;
   16354: out<=1;
   16355: out<=1;
   16356: out<=0;
   16357: out<=1;
   16358: out<=1;
   16359: out<=0;
   16360: out<=1;
   16361: out<=0;
   16362: out<=1;
   16363: out<=0;
   16364: out<=0;
   16365: out<=0;
   16366: out<=1;
   16367: out<=1;
   16368: out<=0;
   16369: out<=1;
   16370: out<=1;
   16371: out<=0;
   16372: out<=0;
   16373: out<=0;
   16374: out<=0;
   16375: out<=0;
   16376: out<=1;
   16377: out<=1;
   16378: out<=0;
   16379: out<=0;
   16380: out<=1;
   16381: out<=0;
   16382: out<=1;
   16383: out<=0;
   16384: out<=1;
   16385: out<=0;
   16386: out<=1;
   16387: out<=0;
   16388: out<=1;
   16389: out<=1;
   16390: out<=0;
   16391: out<=0;
   16392: out<=1;
   16393: out<=1;
   16394: out<=1;
   16395: out<=1;
   16396: out<=1;
   16397: out<=0;
   16398: out<=0;
   16399: out<=1;
   16400: out<=0;
   16401: out<=0;
   16402: out<=1;
   16403: out<=1;
   16404: out<=1;
   16405: out<=0;
   16406: out<=1;
   16407: out<=0;
   16408: out<=1;
   16409: out<=0;
   16410: out<=0;
   16411: out<=1;
   16412: out<=0;
   16413: out<=0;
   16414: out<=0;
   16415: out<=0;
   16416: out<=1;
   16417: out<=1;
   16418: out<=1;
   16419: out<=1;
   16420: out<=0;
   16421: out<=1;
   16422: out<=1;
   16423: out<=0;
   16424: out<=1;
   16425: out<=0;
   16426: out<=1;
   16427: out<=0;
   16428: out<=0;
   16429: out<=0;
   16430: out<=1;
   16431: out<=1;
   16432: out<=0;
   16433: out<=1;
   16434: out<=1;
   16435: out<=0;
   16436: out<=0;
   16437: out<=0;
   16438: out<=0;
   16439: out<=0;
   16440: out<=1;
   16441: out<=1;
   16442: out<=0;
   16443: out<=0;
   16444: out<=1;
   16445: out<=0;
   16446: out<=1;
   16447: out<=0;
   16448: out<=1;
   16449: out<=0;
   16450: out<=1;
   16451: out<=0;
   16452: out<=1;
   16453: out<=1;
   16454: out<=0;
   16455: out<=0;
   16456: out<=1;
   16457: out<=1;
   16458: out<=1;
   16459: out<=1;
   16460: out<=1;
   16461: out<=0;
   16462: out<=0;
   16463: out<=1;
   16464: out<=1;
   16465: out<=1;
   16466: out<=0;
   16467: out<=0;
   16468: out<=0;
   16469: out<=1;
   16470: out<=0;
   16471: out<=1;
   16472: out<=0;
   16473: out<=1;
   16474: out<=1;
   16475: out<=0;
   16476: out<=1;
   16477: out<=1;
   16478: out<=1;
   16479: out<=1;
   16480: out<=0;
   16481: out<=0;
   16482: out<=0;
   16483: out<=0;
   16484: out<=1;
   16485: out<=0;
   16486: out<=0;
   16487: out<=1;
   16488: out<=0;
   16489: out<=1;
   16490: out<=0;
   16491: out<=1;
   16492: out<=1;
   16493: out<=1;
   16494: out<=0;
   16495: out<=0;
   16496: out<=0;
   16497: out<=1;
   16498: out<=1;
   16499: out<=0;
   16500: out<=0;
   16501: out<=0;
   16502: out<=0;
   16503: out<=0;
   16504: out<=1;
   16505: out<=1;
   16506: out<=0;
   16507: out<=0;
   16508: out<=1;
   16509: out<=0;
   16510: out<=1;
   16511: out<=0;
   16512: out<=0;
   16513: out<=1;
   16514: out<=0;
   16515: out<=1;
   16516: out<=0;
   16517: out<=0;
   16518: out<=1;
   16519: out<=1;
   16520: out<=0;
   16521: out<=0;
   16522: out<=0;
   16523: out<=0;
   16524: out<=0;
   16525: out<=1;
   16526: out<=1;
   16527: out<=0;
   16528: out<=0;
   16529: out<=0;
   16530: out<=1;
   16531: out<=1;
   16532: out<=1;
   16533: out<=0;
   16534: out<=1;
   16535: out<=0;
   16536: out<=1;
   16537: out<=0;
   16538: out<=0;
   16539: out<=1;
   16540: out<=0;
   16541: out<=0;
   16542: out<=0;
   16543: out<=0;
   16544: out<=0;
   16545: out<=0;
   16546: out<=0;
   16547: out<=0;
   16548: out<=1;
   16549: out<=0;
   16550: out<=0;
   16551: out<=1;
   16552: out<=0;
   16553: out<=1;
   16554: out<=0;
   16555: out<=1;
   16556: out<=1;
   16557: out<=1;
   16558: out<=0;
   16559: out<=0;
   16560: out<=0;
   16561: out<=1;
   16562: out<=1;
   16563: out<=0;
   16564: out<=0;
   16565: out<=0;
   16566: out<=0;
   16567: out<=0;
   16568: out<=1;
   16569: out<=1;
   16570: out<=0;
   16571: out<=0;
   16572: out<=1;
   16573: out<=0;
   16574: out<=1;
   16575: out<=0;
   16576: out<=0;
   16577: out<=1;
   16578: out<=0;
   16579: out<=1;
   16580: out<=0;
   16581: out<=0;
   16582: out<=1;
   16583: out<=1;
   16584: out<=0;
   16585: out<=0;
   16586: out<=0;
   16587: out<=0;
   16588: out<=0;
   16589: out<=1;
   16590: out<=1;
   16591: out<=0;
   16592: out<=1;
   16593: out<=1;
   16594: out<=0;
   16595: out<=0;
   16596: out<=0;
   16597: out<=1;
   16598: out<=0;
   16599: out<=1;
   16600: out<=0;
   16601: out<=1;
   16602: out<=1;
   16603: out<=0;
   16604: out<=1;
   16605: out<=1;
   16606: out<=1;
   16607: out<=1;
   16608: out<=1;
   16609: out<=1;
   16610: out<=1;
   16611: out<=1;
   16612: out<=0;
   16613: out<=1;
   16614: out<=1;
   16615: out<=0;
   16616: out<=1;
   16617: out<=0;
   16618: out<=1;
   16619: out<=0;
   16620: out<=0;
   16621: out<=0;
   16622: out<=1;
   16623: out<=1;
   16624: out<=0;
   16625: out<=1;
   16626: out<=1;
   16627: out<=0;
   16628: out<=0;
   16629: out<=0;
   16630: out<=0;
   16631: out<=0;
   16632: out<=1;
   16633: out<=1;
   16634: out<=0;
   16635: out<=0;
   16636: out<=1;
   16637: out<=0;
   16638: out<=1;
   16639: out<=0;
   16640: out<=1;
   16641: out<=1;
   16642: out<=0;
   16643: out<=0;
   16644: out<=0;
   16645: out<=1;
   16646: out<=0;
   16647: out<=1;
   16648: out<=0;
   16649: out<=1;
   16650: out<=1;
   16651: out<=0;
   16652: out<=1;
   16653: out<=1;
   16654: out<=1;
   16655: out<=1;
   16656: out<=1;
   16657: out<=0;
   16658: out<=1;
   16659: out<=0;
   16660: out<=1;
   16661: out<=1;
   16662: out<=0;
   16663: out<=0;
   16664: out<=1;
   16665: out<=1;
   16666: out<=1;
   16667: out<=1;
   16668: out<=1;
   16669: out<=0;
   16670: out<=0;
   16671: out<=1;
   16672: out<=0;
   16673: out<=1;
   16674: out<=1;
   16675: out<=0;
   16676: out<=0;
   16677: out<=0;
   16678: out<=0;
   16679: out<=0;
   16680: out<=1;
   16681: out<=1;
   16682: out<=0;
   16683: out<=0;
   16684: out<=1;
   16685: out<=0;
   16686: out<=1;
   16687: out<=0;
   16688: out<=0;
   16689: out<=0;
   16690: out<=0;
   16691: out<=0;
   16692: out<=1;
   16693: out<=0;
   16694: out<=0;
   16695: out<=1;
   16696: out<=0;
   16697: out<=1;
   16698: out<=0;
   16699: out<=1;
   16700: out<=1;
   16701: out<=1;
   16702: out<=0;
   16703: out<=0;
   16704: out<=0;
   16705: out<=0;
   16706: out<=1;
   16707: out<=1;
   16708: out<=1;
   16709: out<=0;
   16710: out<=1;
   16711: out<=0;
   16712: out<=1;
   16713: out<=0;
   16714: out<=0;
   16715: out<=1;
   16716: out<=0;
   16717: out<=0;
   16718: out<=0;
   16719: out<=0;
   16720: out<=1;
   16721: out<=0;
   16722: out<=1;
   16723: out<=0;
   16724: out<=1;
   16725: out<=1;
   16726: out<=0;
   16727: out<=0;
   16728: out<=1;
   16729: out<=1;
   16730: out<=1;
   16731: out<=1;
   16732: out<=1;
   16733: out<=0;
   16734: out<=0;
   16735: out<=1;
   16736: out<=0;
   16737: out<=1;
   16738: out<=1;
   16739: out<=0;
   16740: out<=0;
   16741: out<=0;
   16742: out<=0;
   16743: out<=0;
   16744: out<=1;
   16745: out<=1;
   16746: out<=0;
   16747: out<=0;
   16748: out<=1;
   16749: out<=0;
   16750: out<=1;
   16751: out<=0;
   16752: out<=1;
   16753: out<=1;
   16754: out<=1;
   16755: out<=1;
   16756: out<=0;
   16757: out<=1;
   16758: out<=1;
   16759: out<=0;
   16760: out<=1;
   16761: out<=0;
   16762: out<=1;
   16763: out<=0;
   16764: out<=0;
   16765: out<=0;
   16766: out<=1;
   16767: out<=1;
   16768: out<=1;
   16769: out<=1;
   16770: out<=0;
   16771: out<=0;
   16772: out<=0;
   16773: out<=1;
   16774: out<=0;
   16775: out<=1;
   16776: out<=0;
   16777: out<=1;
   16778: out<=1;
   16779: out<=0;
   16780: out<=1;
   16781: out<=1;
   16782: out<=1;
   16783: out<=1;
   16784: out<=0;
   16785: out<=1;
   16786: out<=0;
   16787: out<=1;
   16788: out<=0;
   16789: out<=0;
   16790: out<=1;
   16791: out<=1;
   16792: out<=0;
   16793: out<=0;
   16794: out<=0;
   16795: out<=0;
   16796: out<=0;
   16797: out<=1;
   16798: out<=1;
   16799: out<=0;
   16800: out<=0;
   16801: out<=1;
   16802: out<=1;
   16803: out<=0;
   16804: out<=0;
   16805: out<=0;
   16806: out<=0;
   16807: out<=0;
   16808: out<=1;
   16809: out<=1;
   16810: out<=0;
   16811: out<=0;
   16812: out<=1;
   16813: out<=0;
   16814: out<=1;
   16815: out<=0;
   16816: out<=1;
   16817: out<=1;
   16818: out<=1;
   16819: out<=1;
   16820: out<=0;
   16821: out<=1;
   16822: out<=1;
   16823: out<=0;
   16824: out<=1;
   16825: out<=0;
   16826: out<=1;
   16827: out<=0;
   16828: out<=0;
   16829: out<=0;
   16830: out<=1;
   16831: out<=1;
   16832: out<=0;
   16833: out<=0;
   16834: out<=1;
   16835: out<=1;
   16836: out<=1;
   16837: out<=0;
   16838: out<=1;
   16839: out<=0;
   16840: out<=1;
   16841: out<=0;
   16842: out<=0;
   16843: out<=1;
   16844: out<=0;
   16845: out<=0;
   16846: out<=0;
   16847: out<=0;
   16848: out<=0;
   16849: out<=1;
   16850: out<=0;
   16851: out<=1;
   16852: out<=0;
   16853: out<=0;
   16854: out<=1;
   16855: out<=1;
   16856: out<=0;
   16857: out<=0;
   16858: out<=0;
   16859: out<=0;
   16860: out<=0;
   16861: out<=1;
   16862: out<=1;
   16863: out<=0;
   16864: out<=0;
   16865: out<=1;
   16866: out<=1;
   16867: out<=0;
   16868: out<=0;
   16869: out<=0;
   16870: out<=0;
   16871: out<=0;
   16872: out<=1;
   16873: out<=1;
   16874: out<=0;
   16875: out<=0;
   16876: out<=1;
   16877: out<=0;
   16878: out<=1;
   16879: out<=0;
   16880: out<=0;
   16881: out<=0;
   16882: out<=0;
   16883: out<=0;
   16884: out<=1;
   16885: out<=0;
   16886: out<=0;
   16887: out<=1;
   16888: out<=0;
   16889: out<=1;
   16890: out<=0;
   16891: out<=1;
   16892: out<=1;
   16893: out<=1;
   16894: out<=0;
   16895: out<=0;
   16896: out<=0;
   16897: out<=0;
   16898: out<=0;
   16899: out<=0;
   16900: out<=1;
   16901: out<=0;
   16902: out<=0;
   16903: out<=1;
   16904: out<=0;
   16905: out<=1;
   16906: out<=0;
   16907: out<=1;
   16908: out<=1;
   16909: out<=1;
   16910: out<=0;
   16911: out<=0;
   16912: out<=0;
   16913: out<=1;
   16914: out<=1;
   16915: out<=0;
   16916: out<=0;
   16917: out<=0;
   16918: out<=0;
   16919: out<=0;
   16920: out<=1;
   16921: out<=1;
   16922: out<=0;
   16923: out<=0;
   16924: out<=1;
   16925: out<=0;
   16926: out<=1;
   16927: out<=0;
   16928: out<=0;
   16929: out<=1;
   16930: out<=0;
   16931: out<=1;
   16932: out<=0;
   16933: out<=0;
   16934: out<=1;
   16935: out<=1;
   16936: out<=0;
   16937: out<=0;
   16938: out<=0;
   16939: out<=0;
   16940: out<=0;
   16941: out<=1;
   16942: out<=1;
   16943: out<=0;
   16944: out<=0;
   16945: out<=0;
   16946: out<=1;
   16947: out<=1;
   16948: out<=1;
   16949: out<=0;
   16950: out<=1;
   16951: out<=0;
   16952: out<=1;
   16953: out<=0;
   16954: out<=0;
   16955: out<=1;
   16956: out<=0;
   16957: out<=0;
   16958: out<=0;
   16959: out<=0;
   16960: out<=1;
   16961: out<=1;
   16962: out<=1;
   16963: out<=1;
   16964: out<=0;
   16965: out<=1;
   16966: out<=1;
   16967: out<=0;
   16968: out<=1;
   16969: out<=0;
   16970: out<=1;
   16971: out<=0;
   16972: out<=0;
   16973: out<=0;
   16974: out<=1;
   16975: out<=1;
   16976: out<=0;
   16977: out<=1;
   16978: out<=1;
   16979: out<=0;
   16980: out<=0;
   16981: out<=0;
   16982: out<=0;
   16983: out<=0;
   16984: out<=1;
   16985: out<=1;
   16986: out<=0;
   16987: out<=0;
   16988: out<=1;
   16989: out<=0;
   16990: out<=1;
   16991: out<=0;
   16992: out<=0;
   16993: out<=1;
   16994: out<=0;
   16995: out<=1;
   16996: out<=0;
   16997: out<=0;
   16998: out<=1;
   16999: out<=1;
   17000: out<=0;
   17001: out<=0;
   17002: out<=0;
   17003: out<=0;
   17004: out<=0;
   17005: out<=1;
   17006: out<=1;
   17007: out<=0;
   17008: out<=1;
   17009: out<=1;
   17010: out<=0;
   17011: out<=0;
   17012: out<=0;
   17013: out<=1;
   17014: out<=0;
   17015: out<=1;
   17016: out<=0;
   17017: out<=1;
   17018: out<=1;
   17019: out<=0;
   17020: out<=1;
   17021: out<=1;
   17022: out<=1;
   17023: out<=1;
   17024: out<=1;
   17025: out<=1;
   17026: out<=1;
   17027: out<=1;
   17028: out<=0;
   17029: out<=1;
   17030: out<=1;
   17031: out<=0;
   17032: out<=1;
   17033: out<=0;
   17034: out<=1;
   17035: out<=0;
   17036: out<=0;
   17037: out<=0;
   17038: out<=1;
   17039: out<=1;
   17040: out<=0;
   17041: out<=1;
   17042: out<=1;
   17043: out<=0;
   17044: out<=0;
   17045: out<=0;
   17046: out<=0;
   17047: out<=0;
   17048: out<=1;
   17049: out<=1;
   17050: out<=0;
   17051: out<=0;
   17052: out<=1;
   17053: out<=0;
   17054: out<=1;
   17055: out<=0;
   17056: out<=1;
   17057: out<=0;
   17058: out<=1;
   17059: out<=0;
   17060: out<=1;
   17061: out<=1;
   17062: out<=0;
   17063: out<=0;
   17064: out<=1;
   17065: out<=1;
   17066: out<=1;
   17067: out<=1;
   17068: out<=1;
   17069: out<=0;
   17070: out<=0;
   17071: out<=1;
   17072: out<=0;
   17073: out<=0;
   17074: out<=1;
   17075: out<=1;
   17076: out<=1;
   17077: out<=0;
   17078: out<=1;
   17079: out<=0;
   17080: out<=1;
   17081: out<=0;
   17082: out<=0;
   17083: out<=1;
   17084: out<=0;
   17085: out<=0;
   17086: out<=0;
   17087: out<=0;
   17088: out<=0;
   17089: out<=0;
   17090: out<=0;
   17091: out<=0;
   17092: out<=1;
   17093: out<=0;
   17094: out<=0;
   17095: out<=1;
   17096: out<=0;
   17097: out<=1;
   17098: out<=0;
   17099: out<=1;
   17100: out<=1;
   17101: out<=1;
   17102: out<=0;
   17103: out<=0;
   17104: out<=0;
   17105: out<=1;
   17106: out<=1;
   17107: out<=0;
   17108: out<=0;
   17109: out<=0;
   17110: out<=0;
   17111: out<=0;
   17112: out<=1;
   17113: out<=1;
   17114: out<=0;
   17115: out<=0;
   17116: out<=1;
   17117: out<=0;
   17118: out<=1;
   17119: out<=0;
   17120: out<=1;
   17121: out<=0;
   17122: out<=1;
   17123: out<=0;
   17124: out<=1;
   17125: out<=1;
   17126: out<=0;
   17127: out<=0;
   17128: out<=1;
   17129: out<=1;
   17130: out<=1;
   17131: out<=1;
   17132: out<=1;
   17133: out<=0;
   17134: out<=0;
   17135: out<=1;
   17136: out<=1;
   17137: out<=1;
   17138: out<=0;
   17139: out<=0;
   17140: out<=0;
   17141: out<=1;
   17142: out<=0;
   17143: out<=1;
   17144: out<=0;
   17145: out<=1;
   17146: out<=1;
   17147: out<=0;
   17148: out<=1;
   17149: out<=1;
   17150: out<=1;
   17151: out<=1;
   17152: out<=0;
   17153: out<=1;
   17154: out<=1;
   17155: out<=0;
   17156: out<=0;
   17157: out<=0;
   17158: out<=0;
   17159: out<=0;
   17160: out<=1;
   17161: out<=1;
   17162: out<=0;
   17163: out<=0;
   17164: out<=1;
   17165: out<=0;
   17166: out<=1;
   17167: out<=0;
   17168: out<=1;
   17169: out<=1;
   17170: out<=1;
   17171: out<=1;
   17172: out<=0;
   17173: out<=1;
   17174: out<=1;
   17175: out<=0;
   17176: out<=1;
   17177: out<=0;
   17178: out<=1;
   17179: out<=0;
   17180: out<=0;
   17181: out<=0;
   17182: out<=1;
   17183: out<=1;
   17184: out<=1;
   17185: out<=1;
   17186: out<=0;
   17187: out<=0;
   17188: out<=0;
   17189: out<=1;
   17190: out<=0;
   17191: out<=1;
   17192: out<=0;
   17193: out<=1;
   17194: out<=1;
   17195: out<=0;
   17196: out<=1;
   17197: out<=1;
   17198: out<=1;
   17199: out<=1;
   17200: out<=0;
   17201: out<=1;
   17202: out<=0;
   17203: out<=1;
   17204: out<=0;
   17205: out<=0;
   17206: out<=1;
   17207: out<=1;
   17208: out<=0;
   17209: out<=0;
   17210: out<=0;
   17211: out<=0;
   17212: out<=0;
   17213: out<=1;
   17214: out<=1;
   17215: out<=0;
   17216: out<=0;
   17217: out<=1;
   17218: out<=1;
   17219: out<=0;
   17220: out<=0;
   17221: out<=0;
   17222: out<=0;
   17223: out<=0;
   17224: out<=1;
   17225: out<=1;
   17226: out<=0;
   17227: out<=0;
   17228: out<=1;
   17229: out<=0;
   17230: out<=1;
   17231: out<=0;
   17232: out<=0;
   17233: out<=0;
   17234: out<=0;
   17235: out<=0;
   17236: out<=1;
   17237: out<=0;
   17238: out<=0;
   17239: out<=1;
   17240: out<=0;
   17241: out<=1;
   17242: out<=0;
   17243: out<=1;
   17244: out<=1;
   17245: out<=1;
   17246: out<=0;
   17247: out<=0;
   17248: out<=0;
   17249: out<=0;
   17250: out<=1;
   17251: out<=1;
   17252: out<=1;
   17253: out<=0;
   17254: out<=1;
   17255: out<=0;
   17256: out<=1;
   17257: out<=0;
   17258: out<=0;
   17259: out<=1;
   17260: out<=0;
   17261: out<=0;
   17262: out<=0;
   17263: out<=0;
   17264: out<=0;
   17265: out<=1;
   17266: out<=0;
   17267: out<=1;
   17268: out<=0;
   17269: out<=0;
   17270: out<=1;
   17271: out<=1;
   17272: out<=0;
   17273: out<=0;
   17274: out<=0;
   17275: out<=0;
   17276: out<=0;
   17277: out<=1;
   17278: out<=1;
   17279: out<=0;
   17280: out<=0;
   17281: out<=1;
   17282: out<=1;
   17283: out<=0;
   17284: out<=0;
   17285: out<=0;
   17286: out<=0;
   17287: out<=0;
   17288: out<=1;
   17289: out<=1;
   17290: out<=0;
   17291: out<=0;
   17292: out<=1;
   17293: out<=0;
   17294: out<=1;
   17295: out<=0;
   17296: out<=0;
   17297: out<=0;
   17298: out<=0;
   17299: out<=0;
   17300: out<=1;
   17301: out<=0;
   17302: out<=0;
   17303: out<=1;
   17304: out<=0;
   17305: out<=1;
   17306: out<=0;
   17307: out<=1;
   17308: out<=1;
   17309: out<=1;
   17310: out<=0;
   17311: out<=0;
   17312: out<=1;
   17313: out<=1;
   17314: out<=0;
   17315: out<=0;
   17316: out<=0;
   17317: out<=1;
   17318: out<=0;
   17319: out<=1;
   17320: out<=0;
   17321: out<=1;
   17322: out<=1;
   17323: out<=0;
   17324: out<=1;
   17325: out<=1;
   17326: out<=1;
   17327: out<=1;
   17328: out<=1;
   17329: out<=0;
   17330: out<=1;
   17331: out<=0;
   17332: out<=1;
   17333: out<=1;
   17334: out<=0;
   17335: out<=0;
   17336: out<=1;
   17337: out<=1;
   17338: out<=1;
   17339: out<=1;
   17340: out<=1;
   17341: out<=0;
   17342: out<=0;
   17343: out<=1;
   17344: out<=0;
   17345: out<=1;
   17346: out<=1;
   17347: out<=0;
   17348: out<=0;
   17349: out<=0;
   17350: out<=0;
   17351: out<=0;
   17352: out<=1;
   17353: out<=1;
   17354: out<=0;
   17355: out<=0;
   17356: out<=1;
   17357: out<=0;
   17358: out<=1;
   17359: out<=0;
   17360: out<=1;
   17361: out<=1;
   17362: out<=1;
   17363: out<=1;
   17364: out<=0;
   17365: out<=1;
   17366: out<=1;
   17367: out<=0;
   17368: out<=1;
   17369: out<=0;
   17370: out<=1;
   17371: out<=0;
   17372: out<=0;
   17373: out<=0;
   17374: out<=1;
   17375: out<=1;
   17376: out<=0;
   17377: out<=0;
   17378: out<=1;
   17379: out<=1;
   17380: out<=1;
   17381: out<=0;
   17382: out<=1;
   17383: out<=0;
   17384: out<=1;
   17385: out<=0;
   17386: out<=0;
   17387: out<=1;
   17388: out<=0;
   17389: out<=0;
   17390: out<=0;
   17391: out<=0;
   17392: out<=1;
   17393: out<=0;
   17394: out<=1;
   17395: out<=0;
   17396: out<=1;
   17397: out<=1;
   17398: out<=0;
   17399: out<=0;
   17400: out<=1;
   17401: out<=1;
   17402: out<=1;
   17403: out<=1;
   17404: out<=1;
   17405: out<=0;
   17406: out<=0;
   17407: out<=1;
   17408: out<=1;
   17409: out<=1;
   17410: out<=0;
   17411: out<=0;
   17412: out<=1;
   17413: out<=0;
   17414: out<=1;
   17415: out<=0;
   17416: out<=1;
   17417: out<=0;
   17418: out<=0;
   17419: out<=1;
   17420: out<=1;
   17421: out<=1;
   17422: out<=1;
   17423: out<=1;
   17424: out<=0;
   17425: out<=1;
   17426: out<=0;
   17427: out<=1;
   17428: out<=1;
   17429: out<=1;
   17430: out<=0;
   17431: out<=0;
   17432: out<=1;
   17433: out<=1;
   17434: out<=1;
   17435: out<=1;
   17436: out<=0;
   17437: out<=1;
   17438: out<=1;
   17439: out<=0;
   17440: out<=1;
   17441: out<=0;
   17442: out<=0;
   17443: out<=1;
   17444: out<=0;
   17445: out<=0;
   17446: out<=0;
   17447: out<=0;
   17448: out<=1;
   17449: out<=1;
   17450: out<=0;
   17451: out<=0;
   17452: out<=0;
   17453: out<=1;
   17454: out<=0;
   17455: out<=1;
   17456: out<=0;
   17457: out<=0;
   17458: out<=0;
   17459: out<=0;
   17460: out<=0;
   17461: out<=1;
   17462: out<=1;
   17463: out<=0;
   17464: out<=1;
   17465: out<=0;
   17466: out<=1;
   17467: out<=0;
   17468: out<=1;
   17469: out<=1;
   17470: out<=0;
   17471: out<=0;
   17472: out<=0;
   17473: out<=0;
   17474: out<=1;
   17475: out<=1;
   17476: out<=0;
   17477: out<=1;
   17478: out<=0;
   17479: out<=1;
   17480: out<=0;
   17481: out<=1;
   17482: out<=1;
   17483: out<=0;
   17484: out<=0;
   17485: out<=0;
   17486: out<=0;
   17487: out<=0;
   17488: out<=0;
   17489: out<=1;
   17490: out<=0;
   17491: out<=1;
   17492: out<=1;
   17493: out<=1;
   17494: out<=0;
   17495: out<=0;
   17496: out<=1;
   17497: out<=1;
   17498: out<=1;
   17499: out<=1;
   17500: out<=0;
   17501: out<=1;
   17502: out<=1;
   17503: out<=0;
   17504: out<=1;
   17505: out<=0;
   17506: out<=0;
   17507: out<=1;
   17508: out<=0;
   17509: out<=0;
   17510: out<=0;
   17511: out<=0;
   17512: out<=1;
   17513: out<=1;
   17514: out<=0;
   17515: out<=0;
   17516: out<=0;
   17517: out<=1;
   17518: out<=0;
   17519: out<=1;
   17520: out<=1;
   17521: out<=1;
   17522: out<=1;
   17523: out<=1;
   17524: out<=1;
   17525: out<=0;
   17526: out<=0;
   17527: out<=1;
   17528: out<=0;
   17529: out<=1;
   17530: out<=0;
   17531: out<=1;
   17532: out<=0;
   17533: out<=0;
   17534: out<=1;
   17535: out<=1;
   17536: out<=1;
   17537: out<=1;
   17538: out<=0;
   17539: out<=0;
   17540: out<=1;
   17541: out<=0;
   17542: out<=1;
   17543: out<=0;
   17544: out<=1;
   17545: out<=0;
   17546: out<=0;
   17547: out<=1;
   17548: out<=1;
   17549: out<=1;
   17550: out<=1;
   17551: out<=1;
   17552: out<=1;
   17553: out<=0;
   17554: out<=1;
   17555: out<=0;
   17556: out<=0;
   17557: out<=0;
   17558: out<=1;
   17559: out<=1;
   17560: out<=0;
   17561: out<=0;
   17562: out<=0;
   17563: out<=0;
   17564: out<=1;
   17565: out<=0;
   17566: out<=0;
   17567: out<=1;
   17568: out<=1;
   17569: out<=0;
   17570: out<=0;
   17571: out<=1;
   17572: out<=0;
   17573: out<=0;
   17574: out<=0;
   17575: out<=0;
   17576: out<=1;
   17577: out<=1;
   17578: out<=0;
   17579: out<=0;
   17580: out<=0;
   17581: out<=1;
   17582: out<=0;
   17583: out<=1;
   17584: out<=1;
   17585: out<=1;
   17586: out<=1;
   17587: out<=1;
   17588: out<=1;
   17589: out<=0;
   17590: out<=0;
   17591: out<=1;
   17592: out<=0;
   17593: out<=1;
   17594: out<=0;
   17595: out<=1;
   17596: out<=0;
   17597: out<=0;
   17598: out<=1;
   17599: out<=1;
   17600: out<=0;
   17601: out<=0;
   17602: out<=1;
   17603: out<=1;
   17604: out<=0;
   17605: out<=1;
   17606: out<=0;
   17607: out<=1;
   17608: out<=0;
   17609: out<=1;
   17610: out<=1;
   17611: out<=0;
   17612: out<=0;
   17613: out<=0;
   17614: out<=0;
   17615: out<=0;
   17616: out<=1;
   17617: out<=0;
   17618: out<=1;
   17619: out<=0;
   17620: out<=0;
   17621: out<=0;
   17622: out<=1;
   17623: out<=1;
   17624: out<=0;
   17625: out<=0;
   17626: out<=0;
   17627: out<=0;
   17628: out<=1;
   17629: out<=0;
   17630: out<=0;
   17631: out<=1;
   17632: out<=1;
   17633: out<=0;
   17634: out<=0;
   17635: out<=1;
   17636: out<=0;
   17637: out<=0;
   17638: out<=0;
   17639: out<=0;
   17640: out<=1;
   17641: out<=1;
   17642: out<=0;
   17643: out<=0;
   17644: out<=0;
   17645: out<=1;
   17646: out<=0;
   17647: out<=1;
   17648: out<=0;
   17649: out<=0;
   17650: out<=0;
   17651: out<=0;
   17652: out<=0;
   17653: out<=1;
   17654: out<=1;
   17655: out<=0;
   17656: out<=1;
   17657: out<=0;
   17658: out<=1;
   17659: out<=0;
   17660: out<=1;
   17661: out<=1;
   17662: out<=0;
   17663: out<=0;
   17664: out<=0;
   17665: out<=1;
   17666: out<=0;
   17667: out<=1;
   17668: out<=1;
   17669: out<=1;
   17670: out<=0;
   17671: out<=0;
   17672: out<=1;
   17673: out<=1;
   17674: out<=1;
   17675: out<=1;
   17676: out<=0;
   17677: out<=1;
   17678: out<=1;
   17679: out<=0;
   17680: out<=0;
   17681: out<=0;
   17682: out<=1;
   17683: out<=1;
   17684: out<=0;
   17685: out<=1;
   17686: out<=0;
   17687: out<=1;
   17688: out<=0;
   17689: out<=1;
   17690: out<=1;
   17691: out<=0;
   17692: out<=0;
   17693: out<=0;
   17694: out<=0;
   17695: out<=0;
   17696: out<=1;
   17697: out<=1;
   17698: out<=1;
   17699: out<=1;
   17700: out<=1;
   17701: out<=0;
   17702: out<=0;
   17703: out<=1;
   17704: out<=0;
   17705: out<=1;
   17706: out<=0;
   17707: out<=1;
   17708: out<=0;
   17709: out<=0;
   17710: out<=1;
   17711: out<=1;
   17712: out<=1;
   17713: out<=0;
   17714: out<=0;
   17715: out<=1;
   17716: out<=0;
   17717: out<=0;
   17718: out<=0;
   17719: out<=0;
   17720: out<=1;
   17721: out<=1;
   17722: out<=0;
   17723: out<=0;
   17724: out<=0;
   17725: out<=1;
   17726: out<=0;
   17727: out<=1;
   17728: out<=0;
   17729: out<=1;
   17730: out<=0;
   17731: out<=1;
   17732: out<=1;
   17733: out<=1;
   17734: out<=0;
   17735: out<=0;
   17736: out<=1;
   17737: out<=1;
   17738: out<=1;
   17739: out<=1;
   17740: out<=0;
   17741: out<=1;
   17742: out<=1;
   17743: out<=0;
   17744: out<=1;
   17745: out<=1;
   17746: out<=0;
   17747: out<=0;
   17748: out<=1;
   17749: out<=0;
   17750: out<=1;
   17751: out<=0;
   17752: out<=1;
   17753: out<=0;
   17754: out<=0;
   17755: out<=1;
   17756: out<=1;
   17757: out<=1;
   17758: out<=1;
   17759: out<=1;
   17760: out<=0;
   17761: out<=0;
   17762: out<=0;
   17763: out<=0;
   17764: out<=0;
   17765: out<=1;
   17766: out<=1;
   17767: out<=0;
   17768: out<=1;
   17769: out<=0;
   17770: out<=1;
   17771: out<=0;
   17772: out<=1;
   17773: out<=1;
   17774: out<=0;
   17775: out<=0;
   17776: out<=1;
   17777: out<=0;
   17778: out<=0;
   17779: out<=1;
   17780: out<=0;
   17781: out<=0;
   17782: out<=0;
   17783: out<=0;
   17784: out<=1;
   17785: out<=1;
   17786: out<=0;
   17787: out<=0;
   17788: out<=0;
   17789: out<=1;
   17790: out<=0;
   17791: out<=1;
   17792: out<=1;
   17793: out<=0;
   17794: out<=1;
   17795: out<=0;
   17796: out<=0;
   17797: out<=0;
   17798: out<=1;
   17799: out<=1;
   17800: out<=0;
   17801: out<=0;
   17802: out<=0;
   17803: out<=0;
   17804: out<=1;
   17805: out<=0;
   17806: out<=0;
   17807: out<=1;
   17808: out<=0;
   17809: out<=0;
   17810: out<=1;
   17811: out<=1;
   17812: out<=0;
   17813: out<=1;
   17814: out<=0;
   17815: out<=1;
   17816: out<=0;
   17817: out<=1;
   17818: out<=1;
   17819: out<=0;
   17820: out<=0;
   17821: out<=0;
   17822: out<=0;
   17823: out<=0;
   17824: out<=0;
   17825: out<=0;
   17826: out<=0;
   17827: out<=0;
   17828: out<=0;
   17829: out<=1;
   17830: out<=1;
   17831: out<=0;
   17832: out<=1;
   17833: out<=0;
   17834: out<=1;
   17835: out<=0;
   17836: out<=1;
   17837: out<=1;
   17838: out<=0;
   17839: out<=0;
   17840: out<=1;
   17841: out<=0;
   17842: out<=0;
   17843: out<=1;
   17844: out<=0;
   17845: out<=0;
   17846: out<=0;
   17847: out<=0;
   17848: out<=1;
   17849: out<=1;
   17850: out<=0;
   17851: out<=0;
   17852: out<=0;
   17853: out<=1;
   17854: out<=0;
   17855: out<=1;
   17856: out<=1;
   17857: out<=0;
   17858: out<=1;
   17859: out<=0;
   17860: out<=0;
   17861: out<=0;
   17862: out<=1;
   17863: out<=1;
   17864: out<=0;
   17865: out<=0;
   17866: out<=0;
   17867: out<=0;
   17868: out<=1;
   17869: out<=0;
   17870: out<=0;
   17871: out<=1;
   17872: out<=1;
   17873: out<=1;
   17874: out<=0;
   17875: out<=0;
   17876: out<=1;
   17877: out<=0;
   17878: out<=1;
   17879: out<=0;
   17880: out<=1;
   17881: out<=0;
   17882: out<=0;
   17883: out<=1;
   17884: out<=1;
   17885: out<=1;
   17886: out<=1;
   17887: out<=1;
   17888: out<=1;
   17889: out<=1;
   17890: out<=1;
   17891: out<=1;
   17892: out<=1;
   17893: out<=0;
   17894: out<=0;
   17895: out<=1;
   17896: out<=0;
   17897: out<=1;
   17898: out<=0;
   17899: out<=1;
   17900: out<=0;
   17901: out<=0;
   17902: out<=1;
   17903: out<=1;
   17904: out<=1;
   17905: out<=0;
   17906: out<=0;
   17907: out<=1;
   17908: out<=0;
   17909: out<=0;
   17910: out<=0;
   17911: out<=0;
   17912: out<=1;
   17913: out<=1;
   17914: out<=0;
   17915: out<=0;
   17916: out<=0;
   17917: out<=1;
   17918: out<=0;
   17919: out<=1;
   17920: out<=1;
   17921: out<=0;
   17922: out<=0;
   17923: out<=1;
   17924: out<=0;
   17925: out<=0;
   17926: out<=0;
   17927: out<=0;
   17928: out<=1;
   17929: out<=1;
   17930: out<=0;
   17931: out<=0;
   17932: out<=0;
   17933: out<=1;
   17934: out<=0;
   17935: out<=1;
   17936: out<=1;
   17937: out<=1;
   17938: out<=1;
   17939: out<=1;
   17940: out<=1;
   17941: out<=0;
   17942: out<=0;
   17943: out<=1;
   17944: out<=0;
   17945: out<=1;
   17946: out<=0;
   17947: out<=1;
   17948: out<=0;
   17949: out<=0;
   17950: out<=1;
   17951: out<=1;
   17952: out<=1;
   17953: out<=1;
   17954: out<=0;
   17955: out<=0;
   17956: out<=1;
   17957: out<=0;
   17958: out<=1;
   17959: out<=0;
   17960: out<=1;
   17961: out<=0;
   17962: out<=0;
   17963: out<=1;
   17964: out<=1;
   17965: out<=1;
   17966: out<=1;
   17967: out<=1;
   17968: out<=1;
   17969: out<=0;
   17970: out<=1;
   17971: out<=0;
   17972: out<=0;
   17973: out<=0;
   17974: out<=1;
   17975: out<=1;
   17976: out<=0;
   17977: out<=0;
   17978: out<=0;
   17979: out<=0;
   17980: out<=1;
   17981: out<=0;
   17982: out<=0;
   17983: out<=1;
   17984: out<=1;
   17985: out<=0;
   17986: out<=0;
   17987: out<=1;
   17988: out<=0;
   17989: out<=0;
   17990: out<=0;
   17991: out<=0;
   17992: out<=1;
   17993: out<=1;
   17994: out<=0;
   17995: out<=0;
   17996: out<=0;
   17997: out<=1;
   17998: out<=0;
   17999: out<=1;
   18000: out<=0;
   18001: out<=0;
   18002: out<=0;
   18003: out<=0;
   18004: out<=0;
   18005: out<=1;
   18006: out<=1;
   18007: out<=0;
   18008: out<=1;
   18009: out<=0;
   18010: out<=1;
   18011: out<=0;
   18012: out<=1;
   18013: out<=1;
   18014: out<=0;
   18015: out<=0;
   18016: out<=0;
   18017: out<=0;
   18018: out<=1;
   18019: out<=1;
   18020: out<=0;
   18021: out<=1;
   18022: out<=0;
   18023: out<=1;
   18024: out<=0;
   18025: out<=1;
   18026: out<=1;
   18027: out<=0;
   18028: out<=0;
   18029: out<=0;
   18030: out<=0;
   18031: out<=0;
   18032: out<=1;
   18033: out<=0;
   18034: out<=1;
   18035: out<=0;
   18036: out<=0;
   18037: out<=0;
   18038: out<=1;
   18039: out<=1;
   18040: out<=0;
   18041: out<=0;
   18042: out<=0;
   18043: out<=0;
   18044: out<=1;
   18045: out<=0;
   18046: out<=0;
   18047: out<=1;
   18048: out<=1;
   18049: out<=0;
   18050: out<=0;
   18051: out<=1;
   18052: out<=0;
   18053: out<=0;
   18054: out<=0;
   18055: out<=0;
   18056: out<=1;
   18057: out<=1;
   18058: out<=0;
   18059: out<=0;
   18060: out<=0;
   18061: out<=1;
   18062: out<=0;
   18063: out<=1;
   18064: out<=0;
   18065: out<=0;
   18066: out<=0;
   18067: out<=0;
   18068: out<=0;
   18069: out<=1;
   18070: out<=1;
   18071: out<=0;
   18072: out<=1;
   18073: out<=0;
   18074: out<=1;
   18075: out<=0;
   18076: out<=1;
   18077: out<=1;
   18078: out<=0;
   18079: out<=0;
   18080: out<=1;
   18081: out<=1;
   18082: out<=0;
   18083: out<=0;
   18084: out<=1;
   18085: out<=0;
   18086: out<=1;
   18087: out<=0;
   18088: out<=1;
   18089: out<=0;
   18090: out<=0;
   18091: out<=1;
   18092: out<=1;
   18093: out<=1;
   18094: out<=1;
   18095: out<=1;
   18096: out<=0;
   18097: out<=1;
   18098: out<=0;
   18099: out<=1;
   18100: out<=1;
   18101: out<=1;
   18102: out<=0;
   18103: out<=0;
   18104: out<=1;
   18105: out<=1;
   18106: out<=1;
   18107: out<=1;
   18108: out<=0;
   18109: out<=1;
   18110: out<=1;
   18111: out<=0;
   18112: out<=1;
   18113: out<=0;
   18114: out<=0;
   18115: out<=1;
   18116: out<=0;
   18117: out<=0;
   18118: out<=0;
   18119: out<=0;
   18120: out<=1;
   18121: out<=1;
   18122: out<=0;
   18123: out<=0;
   18124: out<=0;
   18125: out<=1;
   18126: out<=0;
   18127: out<=1;
   18128: out<=1;
   18129: out<=1;
   18130: out<=1;
   18131: out<=1;
   18132: out<=1;
   18133: out<=0;
   18134: out<=0;
   18135: out<=1;
   18136: out<=0;
   18137: out<=1;
   18138: out<=0;
   18139: out<=1;
   18140: out<=0;
   18141: out<=0;
   18142: out<=1;
   18143: out<=1;
   18144: out<=0;
   18145: out<=0;
   18146: out<=1;
   18147: out<=1;
   18148: out<=0;
   18149: out<=1;
   18150: out<=0;
   18151: out<=1;
   18152: out<=0;
   18153: out<=1;
   18154: out<=1;
   18155: out<=0;
   18156: out<=0;
   18157: out<=0;
   18158: out<=0;
   18159: out<=0;
   18160: out<=0;
   18161: out<=1;
   18162: out<=0;
   18163: out<=1;
   18164: out<=1;
   18165: out<=1;
   18166: out<=0;
   18167: out<=0;
   18168: out<=1;
   18169: out<=1;
   18170: out<=1;
   18171: out<=1;
   18172: out<=0;
   18173: out<=1;
   18174: out<=1;
   18175: out<=0;
   18176: out<=0;
   18177: out<=0;
   18178: out<=0;
   18179: out<=0;
   18180: out<=0;
   18181: out<=1;
   18182: out<=1;
   18183: out<=0;
   18184: out<=1;
   18185: out<=0;
   18186: out<=1;
   18187: out<=0;
   18188: out<=1;
   18189: out<=1;
   18190: out<=0;
   18191: out<=0;
   18192: out<=1;
   18193: out<=0;
   18194: out<=0;
   18195: out<=1;
   18196: out<=0;
   18197: out<=0;
   18198: out<=0;
   18199: out<=0;
   18200: out<=1;
   18201: out<=1;
   18202: out<=0;
   18203: out<=0;
   18204: out<=0;
   18205: out<=1;
   18206: out<=0;
   18207: out<=1;
   18208: out<=1;
   18209: out<=0;
   18210: out<=1;
   18211: out<=0;
   18212: out<=0;
   18213: out<=0;
   18214: out<=1;
   18215: out<=1;
   18216: out<=0;
   18217: out<=0;
   18218: out<=0;
   18219: out<=0;
   18220: out<=1;
   18221: out<=0;
   18222: out<=0;
   18223: out<=1;
   18224: out<=0;
   18225: out<=0;
   18226: out<=1;
   18227: out<=1;
   18228: out<=0;
   18229: out<=1;
   18230: out<=0;
   18231: out<=1;
   18232: out<=0;
   18233: out<=1;
   18234: out<=1;
   18235: out<=0;
   18236: out<=0;
   18237: out<=0;
   18238: out<=0;
   18239: out<=0;
   18240: out<=1;
   18241: out<=1;
   18242: out<=1;
   18243: out<=1;
   18244: out<=1;
   18245: out<=0;
   18246: out<=0;
   18247: out<=1;
   18248: out<=0;
   18249: out<=1;
   18250: out<=0;
   18251: out<=1;
   18252: out<=0;
   18253: out<=0;
   18254: out<=1;
   18255: out<=1;
   18256: out<=1;
   18257: out<=0;
   18258: out<=0;
   18259: out<=1;
   18260: out<=0;
   18261: out<=0;
   18262: out<=0;
   18263: out<=0;
   18264: out<=1;
   18265: out<=1;
   18266: out<=0;
   18267: out<=0;
   18268: out<=0;
   18269: out<=1;
   18270: out<=0;
   18271: out<=1;
   18272: out<=1;
   18273: out<=0;
   18274: out<=1;
   18275: out<=0;
   18276: out<=0;
   18277: out<=0;
   18278: out<=1;
   18279: out<=1;
   18280: out<=0;
   18281: out<=0;
   18282: out<=0;
   18283: out<=0;
   18284: out<=1;
   18285: out<=0;
   18286: out<=0;
   18287: out<=1;
   18288: out<=1;
   18289: out<=1;
   18290: out<=0;
   18291: out<=0;
   18292: out<=1;
   18293: out<=0;
   18294: out<=1;
   18295: out<=0;
   18296: out<=1;
   18297: out<=0;
   18298: out<=0;
   18299: out<=1;
   18300: out<=1;
   18301: out<=1;
   18302: out<=1;
   18303: out<=1;
   18304: out<=1;
   18305: out<=1;
   18306: out<=1;
   18307: out<=1;
   18308: out<=1;
   18309: out<=0;
   18310: out<=0;
   18311: out<=1;
   18312: out<=0;
   18313: out<=1;
   18314: out<=0;
   18315: out<=1;
   18316: out<=0;
   18317: out<=0;
   18318: out<=1;
   18319: out<=1;
   18320: out<=1;
   18321: out<=0;
   18322: out<=0;
   18323: out<=1;
   18324: out<=0;
   18325: out<=0;
   18326: out<=0;
   18327: out<=0;
   18328: out<=1;
   18329: out<=1;
   18330: out<=0;
   18331: out<=0;
   18332: out<=0;
   18333: out<=1;
   18334: out<=0;
   18335: out<=1;
   18336: out<=0;
   18337: out<=1;
   18338: out<=0;
   18339: out<=1;
   18340: out<=1;
   18341: out<=1;
   18342: out<=0;
   18343: out<=0;
   18344: out<=1;
   18345: out<=1;
   18346: out<=1;
   18347: out<=1;
   18348: out<=0;
   18349: out<=1;
   18350: out<=1;
   18351: out<=0;
   18352: out<=0;
   18353: out<=0;
   18354: out<=1;
   18355: out<=1;
   18356: out<=0;
   18357: out<=1;
   18358: out<=0;
   18359: out<=1;
   18360: out<=0;
   18361: out<=1;
   18362: out<=1;
   18363: out<=0;
   18364: out<=0;
   18365: out<=0;
   18366: out<=0;
   18367: out<=0;
   18368: out<=0;
   18369: out<=0;
   18370: out<=0;
   18371: out<=0;
   18372: out<=0;
   18373: out<=1;
   18374: out<=1;
   18375: out<=0;
   18376: out<=1;
   18377: out<=0;
   18378: out<=1;
   18379: out<=0;
   18380: out<=1;
   18381: out<=1;
   18382: out<=0;
   18383: out<=0;
   18384: out<=1;
   18385: out<=0;
   18386: out<=0;
   18387: out<=1;
   18388: out<=0;
   18389: out<=0;
   18390: out<=0;
   18391: out<=0;
   18392: out<=1;
   18393: out<=1;
   18394: out<=0;
   18395: out<=0;
   18396: out<=0;
   18397: out<=1;
   18398: out<=0;
   18399: out<=1;
   18400: out<=0;
   18401: out<=1;
   18402: out<=0;
   18403: out<=1;
   18404: out<=1;
   18405: out<=1;
   18406: out<=0;
   18407: out<=0;
   18408: out<=1;
   18409: out<=1;
   18410: out<=1;
   18411: out<=1;
   18412: out<=0;
   18413: out<=1;
   18414: out<=1;
   18415: out<=0;
   18416: out<=1;
   18417: out<=1;
   18418: out<=0;
   18419: out<=0;
   18420: out<=1;
   18421: out<=0;
   18422: out<=1;
   18423: out<=0;
   18424: out<=1;
   18425: out<=0;
   18426: out<=0;
   18427: out<=1;
   18428: out<=1;
   18429: out<=1;
   18430: out<=1;
   18431: out<=1;
   18432: out<=0;
   18433: out<=0;
   18434: out<=0;
   18435: out<=0;
   18436: out<=0;
   18437: out<=1;
   18438: out<=1;
   18439: out<=0;
   18440: out<=0;
   18441: out<=1;
   18442: out<=0;
   18443: out<=1;
   18444: out<=0;
   18445: out<=0;
   18446: out<=1;
   18447: out<=1;
   18448: out<=1;
   18449: out<=0;
   18450: out<=0;
   18451: out<=1;
   18452: out<=0;
   18453: out<=0;
   18454: out<=0;
   18455: out<=0;
   18456: out<=0;
   18457: out<=0;
   18458: out<=1;
   18459: out<=1;
   18460: out<=1;
   18461: out<=0;
   18462: out<=1;
   18463: out<=0;
   18464: out<=0;
   18465: out<=1;
   18466: out<=0;
   18467: out<=1;
   18468: out<=1;
   18469: out<=1;
   18470: out<=0;
   18471: out<=0;
   18472: out<=0;
   18473: out<=0;
   18474: out<=0;
   18475: out<=0;
   18476: out<=1;
   18477: out<=0;
   18478: out<=0;
   18479: out<=1;
   18480: out<=1;
   18481: out<=1;
   18482: out<=0;
   18483: out<=0;
   18484: out<=1;
   18485: out<=0;
   18486: out<=1;
   18487: out<=0;
   18488: out<=0;
   18489: out<=1;
   18490: out<=1;
   18491: out<=0;
   18492: out<=0;
   18493: out<=0;
   18494: out<=0;
   18495: out<=0;
   18496: out<=1;
   18497: out<=1;
   18498: out<=1;
   18499: out<=1;
   18500: out<=1;
   18501: out<=0;
   18502: out<=0;
   18503: out<=1;
   18504: out<=1;
   18505: out<=0;
   18506: out<=1;
   18507: out<=0;
   18508: out<=1;
   18509: out<=1;
   18510: out<=0;
   18511: out<=0;
   18512: out<=1;
   18513: out<=0;
   18514: out<=0;
   18515: out<=1;
   18516: out<=0;
   18517: out<=0;
   18518: out<=0;
   18519: out<=0;
   18520: out<=0;
   18521: out<=0;
   18522: out<=1;
   18523: out<=1;
   18524: out<=1;
   18525: out<=0;
   18526: out<=1;
   18527: out<=0;
   18528: out<=0;
   18529: out<=1;
   18530: out<=0;
   18531: out<=1;
   18532: out<=1;
   18533: out<=1;
   18534: out<=0;
   18535: out<=0;
   18536: out<=0;
   18537: out<=0;
   18538: out<=0;
   18539: out<=0;
   18540: out<=1;
   18541: out<=0;
   18542: out<=0;
   18543: out<=1;
   18544: out<=0;
   18545: out<=0;
   18546: out<=1;
   18547: out<=1;
   18548: out<=0;
   18549: out<=1;
   18550: out<=0;
   18551: out<=1;
   18552: out<=1;
   18553: out<=0;
   18554: out<=0;
   18555: out<=1;
   18556: out<=1;
   18557: out<=1;
   18558: out<=1;
   18559: out<=1;
   18560: out<=1;
   18561: out<=1;
   18562: out<=1;
   18563: out<=1;
   18564: out<=1;
   18565: out<=0;
   18566: out<=0;
   18567: out<=1;
   18568: out<=1;
   18569: out<=0;
   18570: out<=1;
   18571: out<=0;
   18572: out<=1;
   18573: out<=1;
   18574: out<=0;
   18575: out<=0;
   18576: out<=1;
   18577: out<=0;
   18578: out<=0;
   18579: out<=1;
   18580: out<=0;
   18581: out<=0;
   18582: out<=0;
   18583: out<=0;
   18584: out<=0;
   18585: out<=0;
   18586: out<=1;
   18587: out<=1;
   18588: out<=1;
   18589: out<=0;
   18590: out<=1;
   18591: out<=0;
   18592: out<=1;
   18593: out<=0;
   18594: out<=1;
   18595: out<=0;
   18596: out<=0;
   18597: out<=0;
   18598: out<=1;
   18599: out<=1;
   18600: out<=1;
   18601: out<=1;
   18602: out<=1;
   18603: out<=1;
   18604: out<=0;
   18605: out<=1;
   18606: out<=1;
   18607: out<=0;
   18608: out<=1;
   18609: out<=1;
   18610: out<=0;
   18611: out<=0;
   18612: out<=1;
   18613: out<=0;
   18614: out<=1;
   18615: out<=0;
   18616: out<=0;
   18617: out<=1;
   18618: out<=1;
   18619: out<=0;
   18620: out<=0;
   18621: out<=0;
   18622: out<=0;
   18623: out<=0;
   18624: out<=0;
   18625: out<=0;
   18626: out<=0;
   18627: out<=0;
   18628: out<=0;
   18629: out<=1;
   18630: out<=1;
   18631: out<=0;
   18632: out<=0;
   18633: out<=1;
   18634: out<=0;
   18635: out<=1;
   18636: out<=0;
   18637: out<=0;
   18638: out<=1;
   18639: out<=1;
   18640: out<=1;
   18641: out<=0;
   18642: out<=0;
   18643: out<=1;
   18644: out<=0;
   18645: out<=0;
   18646: out<=0;
   18647: out<=0;
   18648: out<=0;
   18649: out<=0;
   18650: out<=1;
   18651: out<=1;
   18652: out<=1;
   18653: out<=0;
   18654: out<=1;
   18655: out<=0;
   18656: out<=1;
   18657: out<=0;
   18658: out<=1;
   18659: out<=0;
   18660: out<=0;
   18661: out<=0;
   18662: out<=1;
   18663: out<=1;
   18664: out<=1;
   18665: out<=1;
   18666: out<=1;
   18667: out<=1;
   18668: out<=0;
   18669: out<=1;
   18670: out<=1;
   18671: out<=0;
   18672: out<=0;
   18673: out<=0;
   18674: out<=1;
   18675: out<=1;
   18676: out<=0;
   18677: out<=1;
   18678: out<=0;
   18679: out<=1;
   18680: out<=1;
   18681: out<=0;
   18682: out<=0;
   18683: out<=1;
   18684: out<=1;
   18685: out<=1;
   18686: out<=1;
   18687: out<=1;
   18688: out<=1;
   18689: out<=0;
   18690: out<=0;
   18691: out<=1;
   18692: out<=0;
   18693: out<=0;
   18694: out<=0;
   18695: out<=0;
   18696: out<=0;
   18697: out<=0;
   18698: out<=1;
   18699: out<=1;
   18700: out<=1;
   18701: out<=0;
   18702: out<=1;
   18703: out<=0;
   18704: out<=1;
   18705: out<=1;
   18706: out<=1;
   18707: out<=1;
   18708: out<=1;
   18709: out<=0;
   18710: out<=0;
   18711: out<=1;
   18712: out<=1;
   18713: out<=0;
   18714: out<=1;
   18715: out<=0;
   18716: out<=1;
   18717: out<=1;
   18718: out<=0;
   18719: out<=0;
   18720: out<=0;
   18721: out<=0;
   18722: out<=1;
   18723: out<=1;
   18724: out<=0;
   18725: out<=1;
   18726: out<=0;
   18727: out<=1;
   18728: out<=1;
   18729: out<=0;
   18730: out<=0;
   18731: out<=1;
   18732: out<=1;
   18733: out<=1;
   18734: out<=1;
   18735: out<=1;
   18736: out<=0;
   18737: out<=1;
   18738: out<=0;
   18739: out<=1;
   18740: out<=1;
   18741: out<=1;
   18742: out<=0;
   18743: out<=0;
   18744: out<=0;
   18745: out<=0;
   18746: out<=0;
   18747: out<=0;
   18748: out<=1;
   18749: out<=0;
   18750: out<=0;
   18751: out<=1;
   18752: out<=1;
   18753: out<=0;
   18754: out<=0;
   18755: out<=1;
   18756: out<=0;
   18757: out<=0;
   18758: out<=0;
   18759: out<=0;
   18760: out<=0;
   18761: out<=0;
   18762: out<=1;
   18763: out<=1;
   18764: out<=1;
   18765: out<=0;
   18766: out<=1;
   18767: out<=0;
   18768: out<=0;
   18769: out<=0;
   18770: out<=0;
   18771: out<=0;
   18772: out<=0;
   18773: out<=1;
   18774: out<=1;
   18775: out<=0;
   18776: out<=0;
   18777: out<=1;
   18778: out<=0;
   18779: out<=1;
   18780: out<=0;
   18781: out<=0;
   18782: out<=1;
   18783: out<=1;
   18784: out<=1;
   18785: out<=1;
   18786: out<=0;
   18787: out<=0;
   18788: out<=1;
   18789: out<=0;
   18790: out<=1;
   18791: out<=0;
   18792: out<=0;
   18793: out<=1;
   18794: out<=1;
   18795: out<=0;
   18796: out<=0;
   18797: out<=0;
   18798: out<=0;
   18799: out<=0;
   18800: out<=0;
   18801: out<=1;
   18802: out<=0;
   18803: out<=1;
   18804: out<=1;
   18805: out<=1;
   18806: out<=0;
   18807: out<=0;
   18808: out<=0;
   18809: out<=0;
   18810: out<=0;
   18811: out<=0;
   18812: out<=1;
   18813: out<=0;
   18814: out<=0;
   18815: out<=1;
   18816: out<=1;
   18817: out<=0;
   18818: out<=0;
   18819: out<=1;
   18820: out<=0;
   18821: out<=0;
   18822: out<=0;
   18823: out<=0;
   18824: out<=0;
   18825: out<=0;
   18826: out<=1;
   18827: out<=1;
   18828: out<=1;
   18829: out<=0;
   18830: out<=1;
   18831: out<=0;
   18832: out<=0;
   18833: out<=0;
   18834: out<=0;
   18835: out<=0;
   18836: out<=0;
   18837: out<=1;
   18838: out<=1;
   18839: out<=0;
   18840: out<=0;
   18841: out<=1;
   18842: out<=0;
   18843: out<=1;
   18844: out<=0;
   18845: out<=0;
   18846: out<=1;
   18847: out<=1;
   18848: out<=0;
   18849: out<=0;
   18850: out<=1;
   18851: out<=1;
   18852: out<=0;
   18853: out<=1;
   18854: out<=0;
   18855: out<=1;
   18856: out<=1;
   18857: out<=0;
   18858: out<=0;
   18859: out<=1;
   18860: out<=1;
   18861: out<=1;
   18862: out<=1;
   18863: out<=1;
   18864: out<=1;
   18865: out<=0;
   18866: out<=1;
   18867: out<=0;
   18868: out<=0;
   18869: out<=0;
   18870: out<=1;
   18871: out<=1;
   18872: out<=1;
   18873: out<=1;
   18874: out<=1;
   18875: out<=1;
   18876: out<=0;
   18877: out<=1;
   18878: out<=1;
   18879: out<=0;
   18880: out<=1;
   18881: out<=0;
   18882: out<=0;
   18883: out<=1;
   18884: out<=0;
   18885: out<=0;
   18886: out<=0;
   18887: out<=0;
   18888: out<=0;
   18889: out<=0;
   18890: out<=1;
   18891: out<=1;
   18892: out<=1;
   18893: out<=0;
   18894: out<=1;
   18895: out<=0;
   18896: out<=1;
   18897: out<=1;
   18898: out<=1;
   18899: out<=1;
   18900: out<=1;
   18901: out<=0;
   18902: out<=0;
   18903: out<=1;
   18904: out<=1;
   18905: out<=0;
   18906: out<=1;
   18907: out<=0;
   18908: out<=1;
   18909: out<=1;
   18910: out<=0;
   18911: out<=0;
   18912: out<=1;
   18913: out<=1;
   18914: out<=0;
   18915: out<=0;
   18916: out<=1;
   18917: out<=0;
   18918: out<=1;
   18919: out<=0;
   18920: out<=0;
   18921: out<=1;
   18922: out<=1;
   18923: out<=0;
   18924: out<=0;
   18925: out<=0;
   18926: out<=0;
   18927: out<=0;
   18928: out<=1;
   18929: out<=0;
   18930: out<=1;
   18931: out<=0;
   18932: out<=0;
   18933: out<=0;
   18934: out<=1;
   18935: out<=1;
   18936: out<=1;
   18937: out<=1;
   18938: out<=1;
   18939: out<=1;
   18940: out<=0;
   18941: out<=1;
   18942: out<=1;
   18943: out<=0;
   18944: out<=1;
   18945: out<=0;
   18946: out<=1;
   18947: out<=0;
   18948: out<=0;
   18949: out<=0;
   18950: out<=1;
   18951: out<=1;
   18952: out<=1;
   18953: out<=1;
   18954: out<=1;
   18955: out<=1;
   18956: out<=0;
   18957: out<=1;
   18958: out<=1;
   18959: out<=0;
   18960: out<=1;
   18961: out<=1;
   18962: out<=0;
   18963: out<=0;
   18964: out<=1;
   18965: out<=0;
   18966: out<=1;
   18967: out<=0;
   18968: out<=0;
   18969: out<=1;
   18970: out<=1;
   18971: out<=0;
   18972: out<=0;
   18973: out<=0;
   18974: out<=0;
   18975: out<=0;
   18976: out<=1;
   18977: out<=1;
   18978: out<=1;
   18979: out<=1;
   18980: out<=1;
   18981: out<=0;
   18982: out<=0;
   18983: out<=1;
   18984: out<=1;
   18985: out<=0;
   18986: out<=1;
   18987: out<=0;
   18988: out<=1;
   18989: out<=1;
   18990: out<=0;
   18991: out<=0;
   18992: out<=1;
   18993: out<=0;
   18994: out<=0;
   18995: out<=1;
   18996: out<=0;
   18997: out<=0;
   18998: out<=0;
   18999: out<=0;
   19000: out<=0;
   19001: out<=0;
   19002: out<=1;
   19003: out<=1;
   19004: out<=1;
   19005: out<=0;
   19006: out<=1;
   19007: out<=0;
   19008: out<=1;
   19009: out<=0;
   19010: out<=1;
   19011: out<=0;
   19012: out<=0;
   19013: out<=0;
   19014: out<=1;
   19015: out<=1;
   19016: out<=1;
   19017: out<=1;
   19018: out<=1;
   19019: out<=1;
   19020: out<=0;
   19021: out<=1;
   19022: out<=1;
   19023: out<=0;
   19024: out<=0;
   19025: out<=0;
   19026: out<=1;
   19027: out<=1;
   19028: out<=0;
   19029: out<=1;
   19030: out<=0;
   19031: out<=1;
   19032: out<=1;
   19033: out<=0;
   19034: out<=0;
   19035: out<=1;
   19036: out<=1;
   19037: out<=1;
   19038: out<=1;
   19039: out<=1;
   19040: out<=0;
   19041: out<=0;
   19042: out<=0;
   19043: out<=0;
   19044: out<=0;
   19045: out<=1;
   19046: out<=1;
   19047: out<=0;
   19048: out<=0;
   19049: out<=1;
   19050: out<=0;
   19051: out<=1;
   19052: out<=0;
   19053: out<=0;
   19054: out<=1;
   19055: out<=1;
   19056: out<=1;
   19057: out<=0;
   19058: out<=0;
   19059: out<=1;
   19060: out<=0;
   19061: out<=0;
   19062: out<=0;
   19063: out<=0;
   19064: out<=0;
   19065: out<=0;
   19066: out<=1;
   19067: out<=1;
   19068: out<=1;
   19069: out<=0;
   19070: out<=1;
   19071: out<=0;
   19072: out<=0;
   19073: out<=1;
   19074: out<=0;
   19075: out<=1;
   19076: out<=1;
   19077: out<=1;
   19078: out<=0;
   19079: out<=0;
   19080: out<=0;
   19081: out<=0;
   19082: out<=0;
   19083: out<=0;
   19084: out<=1;
   19085: out<=0;
   19086: out<=0;
   19087: out<=1;
   19088: out<=1;
   19089: out<=1;
   19090: out<=0;
   19091: out<=0;
   19092: out<=1;
   19093: out<=0;
   19094: out<=1;
   19095: out<=0;
   19096: out<=0;
   19097: out<=1;
   19098: out<=1;
   19099: out<=0;
   19100: out<=0;
   19101: out<=0;
   19102: out<=0;
   19103: out<=0;
   19104: out<=0;
   19105: out<=0;
   19106: out<=0;
   19107: out<=0;
   19108: out<=0;
   19109: out<=1;
   19110: out<=1;
   19111: out<=0;
   19112: out<=0;
   19113: out<=1;
   19114: out<=0;
   19115: out<=1;
   19116: out<=0;
   19117: out<=0;
   19118: out<=1;
   19119: out<=1;
   19120: out<=1;
   19121: out<=0;
   19122: out<=0;
   19123: out<=1;
   19124: out<=0;
   19125: out<=0;
   19126: out<=0;
   19127: out<=0;
   19128: out<=0;
   19129: out<=0;
   19130: out<=1;
   19131: out<=1;
   19132: out<=1;
   19133: out<=0;
   19134: out<=1;
   19135: out<=0;
   19136: out<=0;
   19137: out<=1;
   19138: out<=0;
   19139: out<=1;
   19140: out<=1;
   19141: out<=1;
   19142: out<=0;
   19143: out<=0;
   19144: out<=0;
   19145: out<=0;
   19146: out<=0;
   19147: out<=0;
   19148: out<=1;
   19149: out<=0;
   19150: out<=0;
   19151: out<=1;
   19152: out<=0;
   19153: out<=0;
   19154: out<=1;
   19155: out<=1;
   19156: out<=0;
   19157: out<=1;
   19158: out<=0;
   19159: out<=1;
   19160: out<=1;
   19161: out<=0;
   19162: out<=0;
   19163: out<=1;
   19164: out<=1;
   19165: out<=1;
   19166: out<=1;
   19167: out<=1;
   19168: out<=1;
   19169: out<=1;
   19170: out<=1;
   19171: out<=1;
   19172: out<=1;
   19173: out<=0;
   19174: out<=0;
   19175: out<=1;
   19176: out<=1;
   19177: out<=0;
   19178: out<=1;
   19179: out<=0;
   19180: out<=1;
   19181: out<=1;
   19182: out<=0;
   19183: out<=0;
   19184: out<=1;
   19185: out<=0;
   19186: out<=0;
   19187: out<=1;
   19188: out<=0;
   19189: out<=0;
   19190: out<=0;
   19191: out<=0;
   19192: out<=0;
   19193: out<=0;
   19194: out<=1;
   19195: out<=1;
   19196: out<=1;
   19197: out<=0;
   19198: out<=1;
   19199: out<=0;
   19200: out<=0;
   19201: out<=0;
   19202: out<=1;
   19203: out<=1;
   19204: out<=0;
   19205: out<=1;
   19206: out<=0;
   19207: out<=1;
   19208: out<=1;
   19209: out<=0;
   19210: out<=0;
   19211: out<=1;
   19212: out<=1;
   19213: out<=1;
   19214: out<=1;
   19215: out<=1;
   19216: out<=1;
   19217: out<=0;
   19218: out<=1;
   19219: out<=0;
   19220: out<=0;
   19221: out<=0;
   19222: out<=1;
   19223: out<=1;
   19224: out<=1;
   19225: out<=1;
   19226: out<=1;
   19227: out<=1;
   19228: out<=0;
   19229: out<=1;
   19230: out<=1;
   19231: out<=0;
   19232: out<=1;
   19233: out<=0;
   19234: out<=0;
   19235: out<=1;
   19236: out<=0;
   19237: out<=0;
   19238: out<=0;
   19239: out<=0;
   19240: out<=0;
   19241: out<=0;
   19242: out<=1;
   19243: out<=1;
   19244: out<=1;
   19245: out<=0;
   19246: out<=1;
   19247: out<=0;
   19248: out<=0;
   19249: out<=0;
   19250: out<=0;
   19251: out<=0;
   19252: out<=0;
   19253: out<=1;
   19254: out<=1;
   19255: out<=0;
   19256: out<=0;
   19257: out<=1;
   19258: out<=0;
   19259: out<=1;
   19260: out<=0;
   19261: out<=0;
   19262: out<=1;
   19263: out<=1;
   19264: out<=1;
   19265: out<=1;
   19266: out<=0;
   19267: out<=0;
   19268: out<=1;
   19269: out<=0;
   19270: out<=1;
   19271: out<=0;
   19272: out<=0;
   19273: out<=1;
   19274: out<=1;
   19275: out<=0;
   19276: out<=0;
   19277: out<=0;
   19278: out<=0;
   19279: out<=0;
   19280: out<=1;
   19281: out<=0;
   19282: out<=1;
   19283: out<=0;
   19284: out<=0;
   19285: out<=0;
   19286: out<=1;
   19287: out<=1;
   19288: out<=1;
   19289: out<=1;
   19290: out<=1;
   19291: out<=1;
   19292: out<=0;
   19293: out<=1;
   19294: out<=1;
   19295: out<=0;
   19296: out<=1;
   19297: out<=0;
   19298: out<=0;
   19299: out<=1;
   19300: out<=0;
   19301: out<=0;
   19302: out<=0;
   19303: out<=0;
   19304: out<=0;
   19305: out<=0;
   19306: out<=1;
   19307: out<=1;
   19308: out<=1;
   19309: out<=0;
   19310: out<=1;
   19311: out<=0;
   19312: out<=1;
   19313: out<=1;
   19314: out<=1;
   19315: out<=1;
   19316: out<=1;
   19317: out<=0;
   19318: out<=0;
   19319: out<=1;
   19320: out<=1;
   19321: out<=0;
   19322: out<=1;
   19323: out<=0;
   19324: out<=1;
   19325: out<=1;
   19326: out<=0;
   19327: out<=0;
   19328: out<=0;
   19329: out<=0;
   19330: out<=1;
   19331: out<=1;
   19332: out<=0;
   19333: out<=1;
   19334: out<=0;
   19335: out<=1;
   19336: out<=1;
   19337: out<=0;
   19338: out<=0;
   19339: out<=1;
   19340: out<=1;
   19341: out<=1;
   19342: out<=1;
   19343: out<=1;
   19344: out<=0;
   19345: out<=1;
   19346: out<=0;
   19347: out<=1;
   19348: out<=1;
   19349: out<=1;
   19350: out<=0;
   19351: out<=0;
   19352: out<=0;
   19353: out<=0;
   19354: out<=0;
   19355: out<=0;
   19356: out<=1;
   19357: out<=0;
   19358: out<=0;
   19359: out<=1;
   19360: out<=1;
   19361: out<=0;
   19362: out<=0;
   19363: out<=1;
   19364: out<=0;
   19365: out<=0;
   19366: out<=0;
   19367: out<=0;
   19368: out<=0;
   19369: out<=0;
   19370: out<=1;
   19371: out<=1;
   19372: out<=1;
   19373: out<=0;
   19374: out<=1;
   19375: out<=0;
   19376: out<=1;
   19377: out<=1;
   19378: out<=1;
   19379: out<=1;
   19380: out<=1;
   19381: out<=0;
   19382: out<=0;
   19383: out<=1;
   19384: out<=1;
   19385: out<=0;
   19386: out<=1;
   19387: out<=0;
   19388: out<=1;
   19389: out<=1;
   19390: out<=0;
   19391: out<=0;
   19392: out<=1;
   19393: out<=1;
   19394: out<=0;
   19395: out<=0;
   19396: out<=1;
   19397: out<=0;
   19398: out<=1;
   19399: out<=0;
   19400: out<=0;
   19401: out<=1;
   19402: out<=1;
   19403: out<=0;
   19404: out<=0;
   19405: out<=0;
   19406: out<=0;
   19407: out<=0;
   19408: out<=0;
   19409: out<=1;
   19410: out<=0;
   19411: out<=1;
   19412: out<=1;
   19413: out<=1;
   19414: out<=0;
   19415: out<=0;
   19416: out<=0;
   19417: out<=0;
   19418: out<=0;
   19419: out<=0;
   19420: out<=1;
   19421: out<=0;
   19422: out<=0;
   19423: out<=1;
   19424: out<=1;
   19425: out<=0;
   19426: out<=0;
   19427: out<=1;
   19428: out<=0;
   19429: out<=0;
   19430: out<=0;
   19431: out<=0;
   19432: out<=0;
   19433: out<=0;
   19434: out<=1;
   19435: out<=1;
   19436: out<=1;
   19437: out<=0;
   19438: out<=1;
   19439: out<=0;
   19440: out<=0;
   19441: out<=0;
   19442: out<=0;
   19443: out<=0;
   19444: out<=0;
   19445: out<=1;
   19446: out<=1;
   19447: out<=0;
   19448: out<=0;
   19449: out<=1;
   19450: out<=0;
   19451: out<=1;
   19452: out<=0;
   19453: out<=0;
   19454: out<=1;
   19455: out<=1;
   19456: out<=0;
   19457: out<=1;
   19458: out<=1;
   19459: out<=0;
   19460: out<=0;
   19461: out<=0;
   19462: out<=0;
   19463: out<=0;
   19464: out<=0;
   19465: out<=0;
   19466: out<=1;
   19467: out<=1;
   19468: out<=0;
   19469: out<=1;
   19470: out<=0;
   19471: out<=1;
   19472: out<=1;
   19473: out<=1;
   19474: out<=1;
   19475: out<=1;
   19476: out<=0;
   19477: out<=1;
   19478: out<=1;
   19479: out<=0;
   19480: out<=0;
   19481: out<=1;
   19482: out<=0;
   19483: out<=1;
   19484: out<=1;
   19485: out<=1;
   19486: out<=0;
   19487: out<=0;
   19488: out<=0;
   19489: out<=0;
   19490: out<=1;
   19491: out<=1;
   19492: out<=1;
   19493: out<=0;
   19494: out<=1;
   19495: out<=0;
   19496: out<=0;
   19497: out<=1;
   19498: out<=1;
   19499: out<=0;
   19500: out<=1;
   19501: out<=1;
   19502: out<=1;
   19503: out<=1;
   19504: out<=1;
   19505: out<=0;
   19506: out<=1;
   19507: out<=0;
   19508: out<=1;
   19509: out<=1;
   19510: out<=0;
   19511: out<=0;
   19512: out<=0;
   19513: out<=0;
   19514: out<=0;
   19515: out<=0;
   19516: out<=0;
   19517: out<=1;
   19518: out<=1;
   19519: out<=0;
   19520: out<=0;
   19521: out<=1;
   19522: out<=1;
   19523: out<=0;
   19524: out<=0;
   19525: out<=0;
   19526: out<=0;
   19527: out<=0;
   19528: out<=0;
   19529: out<=0;
   19530: out<=1;
   19531: out<=1;
   19532: out<=0;
   19533: out<=1;
   19534: out<=0;
   19535: out<=1;
   19536: out<=0;
   19537: out<=0;
   19538: out<=0;
   19539: out<=0;
   19540: out<=1;
   19541: out<=0;
   19542: out<=0;
   19543: out<=1;
   19544: out<=1;
   19545: out<=0;
   19546: out<=1;
   19547: out<=0;
   19548: out<=0;
   19549: out<=0;
   19550: out<=1;
   19551: out<=1;
   19552: out<=1;
   19553: out<=1;
   19554: out<=0;
   19555: out<=0;
   19556: out<=0;
   19557: out<=1;
   19558: out<=0;
   19559: out<=1;
   19560: out<=1;
   19561: out<=0;
   19562: out<=0;
   19563: out<=1;
   19564: out<=0;
   19565: out<=0;
   19566: out<=0;
   19567: out<=0;
   19568: out<=1;
   19569: out<=0;
   19570: out<=1;
   19571: out<=0;
   19572: out<=1;
   19573: out<=1;
   19574: out<=0;
   19575: out<=0;
   19576: out<=0;
   19577: out<=0;
   19578: out<=0;
   19579: out<=0;
   19580: out<=0;
   19581: out<=1;
   19582: out<=1;
   19583: out<=0;
   19584: out<=0;
   19585: out<=1;
   19586: out<=1;
   19587: out<=0;
   19588: out<=0;
   19589: out<=0;
   19590: out<=0;
   19591: out<=0;
   19592: out<=0;
   19593: out<=0;
   19594: out<=1;
   19595: out<=1;
   19596: out<=0;
   19597: out<=1;
   19598: out<=0;
   19599: out<=1;
   19600: out<=0;
   19601: out<=0;
   19602: out<=0;
   19603: out<=0;
   19604: out<=1;
   19605: out<=0;
   19606: out<=0;
   19607: out<=1;
   19608: out<=1;
   19609: out<=0;
   19610: out<=1;
   19611: out<=0;
   19612: out<=0;
   19613: out<=0;
   19614: out<=1;
   19615: out<=1;
   19616: out<=0;
   19617: out<=0;
   19618: out<=1;
   19619: out<=1;
   19620: out<=1;
   19621: out<=0;
   19622: out<=1;
   19623: out<=0;
   19624: out<=0;
   19625: out<=1;
   19626: out<=1;
   19627: out<=0;
   19628: out<=1;
   19629: out<=1;
   19630: out<=1;
   19631: out<=1;
   19632: out<=0;
   19633: out<=1;
   19634: out<=0;
   19635: out<=1;
   19636: out<=0;
   19637: out<=0;
   19638: out<=1;
   19639: out<=1;
   19640: out<=1;
   19641: out<=1;
   19642: out<=1;
   19643: out<=1;
   19644: out<=1;
   19645: out<=0;
   19646: out<=0;
   19647: out<=1;
   19648: out<=0;
   19649: out<=1;
   19650: out<=1;
   19651: out<=0;
   19652: out<=0;
   19653: out<=0;
   19654: out<=0;
   19655: out<=0;
   19656: out<=0;
   19657: out<=0;
   19658: out<=1;
   19659: out<=1;
   19660: out<=0;
   19661: out<=1;
   19662: out<=0;
   19663: out<=1;
   19664: out<=1;
   19665: out<=1;
   19666: out<=1;
   19667: out<=1;
   19668: out<=0;
   19669: out<=1;
   19670: out<=1;
   19671: out<=0;
   19672: out<=0;
   19673: out<=1;
   19674: out<=0;
   19675: out<=1;
   19676: out<=1;
   19677: out<=1;
   19678: out<=0;
   19679: out<=0;
   19680: out<=1;
   19681: out<=1;
   19682: out<=0;
   19683: out<=0;
   19684: out<=0;
   19685: out<=1;
   19686: out<=0;
   19687: out<=1;
   19688: out<=1;
   19689: out<=0;
   19690: out<=0;
   19691: out<=1;
   19692: out<=0;
   19693: out<=0;
   19694: out<=0;
   19695: out<=0;
   19696: out<=0;
   19697: out<=1;
   19698: out<=0;
   19699: out<=1;
   19700: out<=0;
   19701: out<=0;
   19702: out<=1;
   19703: out<=1;
   19704: out<=1;
   19705: out<=1;
   19706: out<=1;
   19707: out<=1;
   19708: out<=1;
   19709: out<=0;
   19710: out<=0;
   19711: out<=1;
   19712: out<=0;
   19713: out<=0;
   19714: out<=0;
   19715: out<=0;
   19716: out<=1;
   19717: out<=0;
   19718: out<=0;
   19719: out<=1;
   19720: out<=1;
   19721: out<=0;
   19722: out<=1;
   19723: out<=0;
   19724: out<=0;
   19725: out<=0;
   19726: out<=1;
   19727: out<=1;
   19728: out<=0;
   19729: out<=1;
   19730: out<=1;
   19731: out<=0;
   19732: out<=0;
   19733: out<=0;
   19734: out<=0;
   19735: out<=0;
   19736: out<=0;
   19737: out<=0;
   19738: out<=1;
   19739: out<=1;
   19740: out<=0;
   19741: out<=1;
   19742: out<=0;
   19743: out<=1;
   19744: out<=1;
   19745: out<=0;
   19746: out<=1;
   19747: out<=0;
   19748: out<=1;
   19749: out<=1;
   19750: out<=0;
   19751: out<=0;
   19752: out<=0;
   19753: out<=0;
   19754: out<=0;
   19755: out<=0;
   19756: out<=0;
   19757: out<=1;
   19758: out<=1;
   19759: out<=0;
   19760: out<=1;
   19761: out<=1;
   19762: out<=0;
   19763: out<=0;
   19764: out<=0;
   19765: out<=1;
   19766: out<=0;
   19767: out<=1;
   19768: out<=1;
   19769: out<=0;
   19770: out<=0;
   19771: out<=1;
   19772: out<=0;
   19773: out<=0;
   19774: out<=0;
   19775: out<=0;
   19776: out<=1;
   19777: out<=1;
   19778: out<=1;
   19779: out<=1;
   19780: out<=0;
   19781: out<=1;
   19782: out<=1;
   19783: out<=0;
   19784: out<=0;
   19785: out<=1;
   19786: out<=0;
   19787: out<=1;
   19788: out<=1;
   19789: out<=1;
   19790: out<=0;
   19791: out<=0;
   19792: out<=0;
   19793: out<=1;
   19794: out<=1;
   19795: out<=0;
   19796: out<=0;
   19797: out<=0;
   19798: out<=0;
   19799: out<=0;
   19800: out<=0;
   19801: out<=0;
   19802: out<=1;
   19803: out<=1;
   19804: out<=0;
   19805: out<=1;
   19806: out<=0;
   19807: out<=1;
   19808: out<=1;
   19809: out<=0;
   19810: out<=1;
   19811: out<=0;
   19812: out<=1;
   19813: out<=1;
   19814: out<=0;
   19815: out<=0;
   19816: out<=0;
   19817: out<=0;
   19818: out<=0;
   19819: out<=0;
   19820: out<=0;
   19821: out<=1;
   19822: out<=1;
   19823: out<=0;
   19824: out<=0;
   19825: out<=0;
   19826: out<=1;
   19827: out<=1;
   19828: out<=1;
   19829: out<=0;
   19830: out<=1;
   19831: out<=0;
   19832: out<=0;
   19833: out<=1;
   19834: out<=1;
   19835: out<=0;
   19836: out<=1;
   19837: out<=1;
   19838: out<=1;
   19839: out<=1;
   19840: out<=1;
   19841: out<=1;
   19842: out<=1;
   19843: out<=1;
   19844: out<=0;
   19845: out<=1;
   19846: out<=1;
   19847: out<=0;
   19848: out<=0;
   19849: out<=1;
   19850: out<=0;
   19851: out<=1;
   19852: out<=1;
   19853: out<=1;
   19854: out<=0;
   19855: out<=0;
   19856: out<=0;
   19857: out<=1;
   19858: out<=1;
   19859: out<=0;
   19860: out<=0;
   19861: out<=0;
   19862: out<=0;
   19863: out<=0;
   19864: out<=0;
   19865: out<=0;
   19866: out<=1;
   19867: out<=1;
   19868: out<=0;
   19869: out<=1;
   19870: out<=0;
   19871: out<=1;
   19872: out<=0;
   19873: out<=1;
   19874: out<=0;
   19875: out<=1;
   19876: out<=0;
   19877: out<=0;
   19878: out<=1;
   19879: out<=1;
   19880: out<=1;
   19881: out<=1;
   19882: out<=1;
   19883: out<=1;
   19884: out<=1;
   19885: out<=0;
   19886: out<=0;
   19887: out<=1;
   19888: out<=1;
   19889: out<=1;
   19890: out<=0;
   19891: out<=0;
   19892: out<=0;
   19893: out<=1;
   19894: out<=0;
   19895: out<=1;
   19896: out<=1;
   19897: out<=0;
   19898: out<=0;
   19899: out<=1;
   19900: out<=0;
   19901: out<=0;
   19902: out<=0;
   19903: out<=0;
   19904: out<=0;
   19905: out<=0;
   19906: out<=0;
   19907: out<=0;
   19908: out<=1;
   19909: out<=0;
   19910: out<=0;
   19911: out<=1;
   19912: out<=1;
   19913: out<=0;
   19914: out<=1;
   19915: out<=0;
   19916: out<=0;
   19917: out<=0;
   19918: out<=1;
   19919: out<=1;
   19920: out<=0;
   19921: out<=1;
   19922: out<=1;
   19923: out<=0;
   19924: out<=0;
   19925: out<=0;
   19926: out<=0;
   19927: out<=0;
   19928: out<=0;
   19929: out<=0;
   19930: out<=1;
   19931: out<=1;
   19932: out<=0;
   19933: out<=1;
   19934: out<=0;
   19935: out<=1;
   19936: out<=0;
   19937: out<=1;
   19938: out<=0;
   19939: out<=1;
   19940: out<=0;
   19941: out<=0;
   19942: out<=1;
   19943: out<=1;
   19944: out<=1;
   19945: out<=1;
   19946: out<=1;
   19947: out<=1;
   19948: out<=1;
   19949: out<=0;
   19950: out<=0;
   19951: out<=1;
   19952: out<=0;
   19953: out<=0;
   19954: out<=1;
   19955: out<=1;
   19956: out<=1;
   19957: out<=0;
   19958: out<=1;
   19959: out<=0;
   19960: out<=0;
   19961: out<=1;
   19962: out<=1;
   19963: out<=0;
   19964: out<=1;
   19965: out<=1;
   19966: out<=1;
   19967: out<=1;
   19968: out<=0;
   19969: out<=0;
   19970: out<=1;
   19971: out<=1;
   19972: out<=1;
   19973: out<=0;
   19974: out<=1;
   19975: out<=0;
   19976: out<=0;
   19977: out<=1;
   19978: out<=1;
   19979: out<=0;
   19980: out<=1;
   19981: out<=1;
   19982: out<=1;
   19983: out<=1;
   19984: out<=0;
   19985: out<=1;
   19986: out<=0;
   19987: out<=1;
   19988: out<=0;
   19989: out<=0;
   19990: out<=1;
   19991: out<=1;
   19992: out<=1;
   19993: out<=1;
   19994: out<=1;
   19995: out<=1;
   19996: out<=1;
   19997: out<=0;
   19998: out<=0;
   19999: out<=1;
   20000: out<=0;
   20001: out<=1;
   20002: out<=1;
   20003: out<=0;
   20004: out<=0;
   20005: out<=0;
   20006: out<=0;
   20007: out<=0;
   20008: out<=0;
   20009: out<=0;
   20010: out<=1;
   20011: out<=1;
   20012: out<=0;
   20013: out<=1;
   20014: out<=0;
   20015: out<=1;
   20016: out<=0;
   20017: out<=0;
   20018: out<=0;
   20019: out<=0;
   20020: out<=1;
   20021: out<=0;
   20022: out<=0;
   20023: out<=1;
   20024: out<=1;
   20025: out<=0;
   20026: out<=1;
   20027: out<=0;
   20028: out<=0;
   20029: out<=0;
   20030: out<=1;
   20031: out<=1;
   20032: out<=1;
   20033: out<=1;
   20034: out<=0;
   20035: out<=0;
   20036: out<=0;
   20037: out<=1;
   20038: out<=0;
   20039: out<=1;
   20040: out<=1;
   20041: out<=0;
   20042: out<=0;
   20043: out<=1;
   20044: out<=0;
   20045: out<=0;
   20046: out<=0;
   20047: out<=0;
   20048: out<=0;
   20049: out<=1;
   20050: out<=0;
   20051: out<=1;
   20052: out<=0;
   20053: out<=0;
   20054: out<=1;
   20055: out<=1;
   20056: out<=1;
   20057: out<=1;
   20058: out<=1;
   20059: out<=1;
   20060: out<=1;
   20061: out<=0;
   20062: out<=0;
   20063: out<=1;
   20064: out<=0;
   20065: out<=1;
   20066: out<=1;
   20067: out<=0;
   20068: out<=0;
   20069: out<=0;
   20070: out<=0;
   20071: out<=0;
   20072: out<=0;
   20073: out<=0;
   20074: out<=1;
   20075: out<=1;
   20076: out<=0;
   20077: out<=1;
   20078: out<=0;
   20079: out<=1;
   20080: out<=1;
   20081: out<=1;
   20082: out<=1;
   20083: out<=1;
   20084: out<=0;
   20085: out<=1;
   20086: out<=1;
   20087: out<=0;
   20088: out<=0;
   20089: out<=1;
   20090: out<=0;
   20091: out<=1;
   20092: out<=1;
   20093: out<=1;
   20094: out<=0;
   20095: out<=0;
   20096: out<=0;
   20097: out<=0;
   20098: out<=1;
   20099: out<=1;
   20100: out<=1;
   20101: out<=0;
   20102: out<=1;
   20103: out<=0;
   20104: out<=0;
   20105: out<=1;
   20106: out<=1;
   20107: out<=0;
   20108: out<=1;
   20109: out<=1;
   20110: out<=1;
   20111: out<=1;
   20112: out<=1;
   20113: out<=0;
   20114: out<=1;
   20115: out<=0;
   20116: out<=1;
   20117: out<=1;
   20118: out<=0;
   20119: out<=0;
   20120: out<=0;
   20121: out<=0;
   20122: out<=0;
   20123: out<=0;
   20124: out<=0;
   20125: out<=1;
   20126: out<=1;
   20127: out<=0;
   20128: out<=0;
   20129: out<=1;
   20130: out<=1;
   20131: out<=0;
   20132: out<=0;
   20133: out<=0;
   20134: out<=0;
   20135: out<=0;
   20136: out<=0;
   20137: out<=0;
   20138: out<=1;
   20139: out<=1;
   20140: out<=0;
   20141: out<=1;
   20142: out<=0;
   20143: out<=1;
   20144: out<=1;
   20145: out<=1;
   20146: out<=1;
   20147: out<=1;
   20148: out<=0;
   20149: out<=1;
   20150: out<=1;
   20151: out<=0;
   20152: out<=0;
   20153: out<=1;
   20154: out<=0;
   20155: out<=1;
   20156: out<=1;
   20157: out<=1;
   20158: out<=0;
   20159: out<=0;
   20160: out<=1;
   20161: out<=1;
   20162: out<=0;
   20163: out<=0;
   20164: out<=0;
   20165: out<=1;
   20166: out<=0;
   20167: out<=1;
   20168: out<=1;
   20169: out<=0;
   20170: out<=0;
   20171: out<=1;
   20172: out<=0;
   20173: out<=0;
   20174: out<=0;
   20175: out<=0;
   20176: out<=1;
   20177: out<=0;
   20178: out<=1;
   20179: out<=0;
   20180: out<=1;
   20181: out<=1;
   20182: out<=0;
   20183: out<=0;
   20184: out<=0;
   20185: out<=0;
   20186: out<=0;
   20187: out<=0;
   20188: out<=0;
   20189: out<=1;
   20190: out<=1;
   20191: out<=0;
   20192: out<=0;
   20193: out<=1;
   20194: out<=1;
   20195: out<=0;
   20196: out<=0;
   20197: out<=0;
   20198: out<=0;
   20199: out<=0;
   20200: out<=0;
   20201: out<=0;
   20202: out<=1;
   20203: out<=1;
   20204: out<=0;
   20205: out<=1;
   20206: out<=0;
   20207: out<=1;
   20208: out<=0;
   20209: out<=0;
   20210: out<=0;
   20211: out<=0;
   20212: out<=1;
   20213: out<=0;
   20214: out<=0;
   20215: out<=1;
   20216: out<=1;
   20217: out<=0;
   20218: out<=1;
   20219: out<=0;
   20220: out<=0;
   20221: out<=0;
   20222: out<=1;
   20223: out<=1;
   20224: out<=0;
   20225: out<=1;
   20226: out<=0;
   20227: out<=1;
   20228: out<=0;
   20229: out<=0;
   20230: out<=1;
   20231: out<=1;
   20232: out<=1;
   20233: out<=1;
   20234: out<=1;
   20235: out<=1;
   20236: out<=1;
   20237: out<=0;
   20238: out<=0;
   20239: out<=1;
   20240: out<=1;
   20241: out<=1;
   20242: out<=0;
   20243: out<=0;
   20244: out<=0;
   20245: out<=1;
   20246: out<=0;
   20247: out<=1;
   20248: out<=1;
   20249: out<=0;
   20250: out<=0;
   20251: out<=1;
   20252: out<=0;
   20253: out<=0;
   20254: out<=0;
   20255: out<=0;
   20256: out<=1;
   20257: out<=1;
   20258: out<=1;
   20259: out<=1;
   20260: out<=0;
   20261: out<=1;
   20262: out<=1;
   20263: out<=0;
   20264: out<=0;
   20265: out<=1;
   20266: out<=0;
   20267: out<=1;
   20268: out<=1;
   20269: out<=1;
   20270: out<=0;
   20271: out<=0;
   20272: out<=0;
   20273: out<=1;
   20274: out<=1;
   20275: out<=0;
   20276: out<=0;
   20277: out<=0;
   20278: out<=0;
   20279: out<=0;
   20280: out<=0;
   20281: out<=0;
   20282: out<=1;
   20283: out<=1;
   20284: out<=0;
   20285: out<=1;
   20286: out<=0;
   20287: out<=1;
   20288: out<=0;
   20289: out<=1;
   20290: out<=0;
   20291: out<=1;
   20292: out<=0;
   20293: out<=0;
   20294: out<=1;
   20295: out<=1;
   20296: out<=1;
   20297: out<=1;
   20298: out<=1;
   20299: out<=1;
   20300: out<=1;
   20301: out<=0;
   20302: out<=0;
   20303: out<=1;
   20304: out<=0;
   20305: out<=0;
   20306: out<=1;
   20307: out<=1;
   20308: out<=1;
   20309: out<=0;
   20310: out<=1;
   20311: out<=0;
   20312: out<=0;
   20313: out<=1;
   20314: out<=1;
   20315: out<=0;
   20316: out<=1;
   20317: out<=1;
   20318: out<=1;
   20319: out<=1;
   20320: out<=0;
   20321: out<=0;
   20322: out<=0;
   20323: out<=0;
   20324: out<=1;
   20325: out<=0;
   20326: out<=0;
   20327: out<=1;
   20328: out<=1;
   20329: out<=0;
   20330: out<=1;
   20331: out<=0;
   20332: out<=0;
   20333: out<=0;
   20334: out<=1;
   20335: out<=1;
   20336: out<=0;
   20337: out<=1;
   20338: out<=1;
   20339: out<=0;
   20340: out<=0;
   20341: out<=0;
   20342: out<=0;
   20343: out<=0;
   20344: out<=0;
   20345: out<=0;
   20346: out<=1;
   20347: out<=1;
   20348: out<=0;
   20349: out<=1;
   20350: out<=0;
   20351: out<=1;
   20352: out<=1;
   20353: out<=0;
   20354: out<=1;
   20355: out<=0;
   20356: out<=1;
   20357: out<=1;
   20358: out<=0;
   20359: out<=0;
   20360: out<=0;
   20361: out<=0;
   20362: out<=0;
   20363: out<=0;
   20364: out<=0;
   20365: out<=1;
   20366: out<=1;
   20367: out<=0;
   20368: out<=1;
   20369: out<=1;
   20370: out<=0;
   20371: out<=0;
   20372: out<=0;
   20373: out<=1;
   20374: out<=0;
   20375: out<=1;
   20376: out<=1;
   20377: out<=0;
   20378: out<=0;
   20379: out<=1;
   20380: out<=0;
   20381: out<=0;
   20382: out<=0;
   20383: out<=0;
   20384: out<=0;
   20385: out<=0;
   20386: out<=0;
   20387: out<=0;
   20388: out<=1;
   20389: out<=0;
   20390: out<=0;
   20391: out<=1;
   20392: out<=1;
   20393: out<=0;
   20394: out<=1;
   20395: out<=0;
   20396: out<=0;
   20397: out<=0;
   20398: out<=1;
   20399: out<=1;
   20400: out<=0;
   20401: out<=1;
   20402: out<=1;
   20403: out<=0;
   20404: out<=0;
   20405: out<=0;
   20406: out<=0;
   20407: out<=0;
   20408: out<=0;
   20409: out<=0;
   20410: out<=1;
   20411: out<=1;
   20412: out<=0;
   20413: out<=1;
   20414: out<=0;
   20415: out<=1;
   20416: out<=1;
   20417: out<=0;
   20418: out<=1;
   20419: out<=0;
   20420: out<=1;
   20421: out<=1;
   20422: out<=0;
   20423: out<=0;
   20424: out<=0;
   20425: out<=0;
   20426: out<=0;
   20427: out<=0;
   20428: out<=0;
   20429: out<=1;
   20430: out<=1;
   20431: out<=0;
   20432: out<=0;
   20433: out<=0;
   20434: out<=1;
   20435: out<=1;
   20436: out<=1;
   20437: out<=0;
   20438: out<=1;
   20439: out<=0;
   20440: out<=0;
   20441: out<=1;
   20442: out<=1;
   20443: out<=0;
   20444: out<=1;
   20445: out<=1;
   20446: out<=1;
   20447: out<=1;
   20448: out<=1;
   20449: out<=1;
   20450: out<=1;
   20451: out<=1;
   20452: out<=0;
   20453: out<=1;
   20454: out<=1;
   20455: out<=0;
   20456: out<=0;
   20457: out<=1;
   20458: out<=0;
   20459: out<=1;
   20460: out<=1;
   20461: out<=1;
   20462: out<=0;
   20463: out<=0;
   20464: out<=0;
   20465: out<=1;
   20466: out<=1;
   20467: out<=0;
   20468: out<=0;
   20469: out<=0;
   20470: out<=0;
   20471: out<=0;
   20472: out<=0;
   20473: out<=0;
   20474: out<=1;
   20475: out<=1;
   20476: out<=0;
   20477: out<=1;
   20478: out<=0;
   20479: out<=1;
   20480: out<=1;
   20481: out<=0;
   20482: out<=1;
   20483: out<=0;
   20484: out<=0;
   20485: out<=0;
   20486: out<=1;
   20487: out<=1;
   20488: out<=0;
   20489: out<=0;
   20490: out<=0;
   20491: out<=0;
   20492: out<=1;
   20493: out<=0;
   20494: out<=0;
   20495: out<=1;
   20496: out<=0;
   20497: out<=0;
   20498: out<=1;
   20499: out<=1;
   20500: out<=0;
   20501: out<=1;
   20502: out<=0;
   20503: out<=1;
   20504: out<=0;
   20505: out<=1;
   20506: out<=1;
   20507: out<=0;
   20508: out<=0;
   20509: out<=0;
   20510: out<=0;
   20511: out<=0;
   20512: out<=1;
   20513: out<=1;
   20514: out<=1;
   20515: out<=1;
   20516: out<=1;
   20517: out<=0;
   20518: out<=0;
   20519: out<=1;
   20520: out<=0;
   20521: out<=1;
   20522: out<=0;
   20523: out<=1;
   20524: out<=0;
   20525: out<=0;
   20526: out<=1;
   20527: out<=1;
   20528: out<=0;
   20529: out<=1;
   20530: out<=1;
   20531: out<=0;
   20532: out<=1;
   20533: out<=1;
   20534: out<=1;
   20535: out<=1;
   20536: out<=0;
   20537: out<=0;
   20538: out<=1;
   20539: out<=1;
   20540: out<=1;
   20541: out<=0;
   20542: out<=1;
   20543: out<=0;
   20544: out<=1;
   20545: out<=0;
   20546: out<=1;
   20547: out<=0;
   20548: out<=0;
   20549: out<=0;
   20550: out<=1;
   20551: out<=1;
   20552: out<=0;
   20553: out<=0;
   20554: out<=0;
   20555: out<=0;
   20556: out<=1;
   20557: out<=0;
   20558: out<=0;
   20559: out<=1;
   20560: out<=1;
   20561: out<=1;
   20562: out<=0;
   20563: out<=0;
   20564: out<=1;
   20565: out<=0;
   20566: out<=1;
   20567: out<=0;
   20568: out<=1;
   20569: out<=0;
   20570: out<=0;
   20571: out<=1;
   20572: out<=1;
   20573: out<=1;
   20574: out<=1;
   20575: out<=1;
   20576: out<=0;
   20577: out<=0;
   20578: out<=0;
   20579: out<=0;
   20580: out<=0;
   20581: out<=1;
   20582: out<=1;
   20583: out<=0;
   20584: out<=1;
   20585: out<=0;
   20586: out<=1;
   20587: out<=0;
   20588: out<=1;
   20589: out<=1;
   20590: out<=0;
   20591: out<=0;
   20592: out<=0;
   20593: out<=1;
   20594: out<=1;
   20595: out<=0;
   20596: out<=1;
   20597: out<=1;
   20598: out<=1;
   20599: out<=1;
   20600: out<=0;
   20601: out<=0;
   20602: out<=1;
   20603: out<=1;
   20604: out<=1;
   20605: out<=0;
   20606: out<=1;
   20607: out<=0;
   20608: out<=0;
   20609: out<=1;
   20610: out<=0;
   20611: out<=1;
   20612: out<=1;
   20613: out<=1;
   20614: out<=0;
   20615: out<=0;
   20616: out<=1;
   20617: out<=1;
   20618: out<=1;
   20619: out<=1;
   20620: out<=0;
   20621: out<=1;
   20622: out<=1;
   20623: out<=0;
   20624: out<=0;
   20625: out<=0;
   20626: out<=1;
   20627: out<=1;
   20628: out<=0;
   20629: out<=1;
   20630: out<=0;
   20631: out<=1;
   20632: out<=0;
   20633: out<=1;
   20634: out<=1;
   20635: out<=0;
   20636: out<=0;
   20637: out<=0;
   20638: out<=0;
   20639: out<=0;
   20640: out<=0;
   20641: out<=0;
   20642: out<=0;
   20643: out<=0;
   20644: out<=0;
   20645: out<=1;
   20646: out<=1;
   20647: out<=0;
   20648: out<=1;
   20649: out<=0;
   20650: out<=1;
   20651: out<=0;
   20652: out<=1;
   20653: out<=1;
   20654: out<=0;
   20655: out<=0;
   20656: out<=0;
   20657: out<=1;
   20658: out<=1;
   20659: out<=0;
   20660: out<=1;
   20661: out<=1;
   20662: out<=1;
   20663: out<=1;
   20664: out<=0;
   20665: out<=0;
   20666: out<=1;
   20667: out<=1;
   20668: out<=1;
   20669: out<=0;
   20670: out<=1;
   20671: out<=0;
   20672: out<=0;
   20673: out<=1;
   20674: out<=0;
   20675: out<=1;
   20676: out<=1;
   20677: out<=1;
   20678: out<=0;
   20679: out<=0;
   20680: out<=1;
   20681: out<=1;
   20682: out<=1;
   20683: out<=1;
   20684: out<=0;
   20685: out<=1;
   20686: out<=1;
   20687: out<=0;
   20688: out<=1;
   20689: out<=1;
   20690: out<=0;
   20691: out<=0;
   20692: out<=1;
   20693: out<=0;
   20694: out<=1;
   20695: out<=0;
   20696: out<=1;
   20697: out<=0;
   20698: out<=0;
   20699: out<=1;
   20700: out<=1;
   20701: out<=1;
   20702: out<=1;
   20703: out<=1;
   20704: out<=1;
   20705: out<=1;
   20706: out<=1;
   20707: out<=1;
   20708: out<=1;
   20709: out<=0;
   20710: out<=0;
   20711: out<=1;
   20712: out<=0;
   20713: out<=1;
   20714: out<=0;
   20715: out<=1;
   20716: out<=0;
   20717: out<=0;
   20718: out<=1;
   20719: out<=1;
   20720: out<=0;
   20721: out<=1;
   20722: out<=1;
   20723: out<=0;
   20724: out<=1;
   20725: out<=1;
   20726: out<=1;
   20727: out<=1;
   20728: out<=0;
   20729: out<=0;
   20730: out<=1;
   20731: out<=1;
   20732: out<=1;
   20733: out<=0;
   20734: out<=1;
   20735: out<=0;
   20736: out<=1;
   20737: out<=1;
   20738: out<=0;
   20739: out<=0;
   20740: out<=1;
   20741: out<=0;
   20742: out<=1;
   20743: out<=0;
   20744: out<=1;
   20745: out<=0;
   20746: out<=0;
   20747: out<=1;
   20748: out<=1;
   20749: out<=1;
   20750: out<=1;
   20751: out<=1;
   20752: out<=1;
   20753: out<=0;
   20754: out<=1;
   20755: out<=0;
   20756: out<=0;
   20757: out<=0;
   20758: out<=1;
   20759: out<=1;
   20760: out<=0;
   20761: out<=0;
   20762: out<=0;
   20763: out<=0;
   20764: out<=1;
   20765: out<=0;
   20766: out<=0;
   20767: out<=1;
   20768: out<=0;
   20769: out<=1;
   20770: out<=1;
   20771: out<=0;
   20772: out<=1;
   20773: out<=1;
   20774: out<=1;
   20775: out<=1;
   20776: out<=0;
   20777: out<=0;
   20778: out<=1;
   20779: out<=1;
   20780: out<=1;
   20781: out<=0;
   20782: out<=1;
   20783: out<=0;
   20784: out<=0;
   20785: out<=0;
   20786: out<=0;
   20787: out<=0;
   20788: out<=0;
   20789: out<=1;
   20790: out<=1;
   20791: out<=0;
   20792: out<=1;
   20793: out<=0;
   20794: out<=1;
   20795: out<=0;
   20796: out<=1;
   20797: out<=1;
   20798: out<=0;
   20799: out<=0;
   20800: out<=0;
   20801: out<=0;
   20802: out<=1;
   20803: out<=1;
   20804: out<=0;
   20805: out<=1;
   20806: out<=0;
   20807: out<=1;
   20808: out<=0;
   20809: out<=1;
   20810: out<=1;
   20811: out<=0;
   20812: out<=0;
   20813: out<=0;
   20814: out<=0;
   20815: out<=0;
   20816: out<=1;
   20817: out<=0;
   20818: out<=1;
   20819: out<=0;
   20820: out<=0;
   20821: out<=0;
   20822: out<=1;
   20823: out<=1;
   20824: out<=0;
   20825: out<=0;
   20826: out<=0;
   20827: out<=0;
   20828: out<=1;
   20829: out<=0;
   20830: out<=0;
   20831: out<=1;
   20832: out<=0;
   20833: out<=1;
   20834: out<=1;
   20835: out<=0;
   20836: out<=1;
   20837: out<=1;
   20838: out<=1;
   20839: out<=1;
   20840: out<=0;
   20841: out<=0;
   20842: out<=1;
   20843: out<=1;
   20844: out<=1;
   20845: out<=0;
   20846: out<=1;
   20847: out<=0;
   20848: out<=1;
   20849: out<=1;
   20850: out<=1;
   20851: out<=1;
   20852: out<=1;
   20853: out<=0;
   20854: out<=0;
   20855: out<=1;
   20856: out<=0;
   20857: out<=1;
   20858: out<=0;
   20859: out<=1;
   20860: out<=0;
   20861: out<=0;
   20862: out<=1;
   20863: out<=1;
   20864: out<=1;
   20865: out<=1;
   20866: out<=0;
   20867: out<=0;
   20868: out<=1;
   20869: out<=0;
   20870: out<=1;
   20871: out<=0;
   20872: out<=1;
   20873: out<=0;
   20874: out<=0;
   20875: out<=1;
   20876: out<=1;
   20877: out<=1;
   20878: out<=1;
   20879: out<=1;
   20880: out<=0;
   20881: out<=1;
   20882: out<=0;
   20883: out<=1;
   20884: out<=1;
   20885: out<=1;
   20886: out<=0;
   20887: out<=0;
   20888: out<=1;
   20889: out<=1;
   20890: out<=1;
   20891: out<=1;
   20892: out<=0;
   20893: out<=1;
   20894: out<=1;
   20895: out<=0;
   20896: out<=0;
   20897: out<=1;
   20898: out<=1;
   20899: out<=0;
   20900: out<=1;
   20901: out<=1;
   20902: out<=1;
   20903: out<=1;
   20904: out<=0;
   20905: out<=0;
   20906: out<=1;
   20907: out<=1;
   20908: out<=1;
   20909: out<=0;
   20910: out<=1;
   20911: out<=0;
   20912: out<=1;
   20913: out<=1;
   20914: out<=1;
   20915: out<=1;
   20916: out<=1;
   20917: out<=0;
   20918: out<=0;
   20919: out<=1;
   20920: out<=0;
   20921: out<=1;
   20922: out<=0;
   20923: out<=1;
   20924: out<=0;
   20925: out<=0;
   20926: out<=1;
   20927: out<=1;
   20928: out<=0;
   20929: out<=0;
   20930: out<=1;
   20931: out<=1;
   20932: out<=0;
   20933: out<=1;
   20934: out<=0;
   20935: out<=1;
   20936: out<=0;
   20937: out<=1;
   20938: out<=1;
   20939: out<=0;
   20940: out<=0;
   20941: out<=0;
   20942: out<=0;
   20943: out<=0;
   20944: out<=0;
   20945: out<=1;
   20946: out<=0;
   20947: out<=1;
   20948: out<=1;
   20949: out<=1;
   20950: out<=0;
   20951: out<=0;
   20952: out<=1;
   20953: out<=1;
   20954: out<=1;
   20955: out<=1;
   20956: out<=0;
   20957: out<=1;
   20958: out<=1;
   20959: out<=0;
   20960: out<=0;
   20961: out<=1;
   20962: out<=1;
   20963: out<=0;
   20964: out<=1;
   20965: out<=1;
   20966: out<=1;
   20967: out<=1;
   20968: out<=0;
   20969: out<=0;
   20970: out<=1;
   20971: out<=1;
   20972: out<=1;
   20973: out<=0;
   20974: out<=1;
   20975: out<=0;
   20976: out<=0;
   20977: out<=0;
   20978: out<=0;
   20979: out<=0;
   20980: out<=0;
   20981: out<=1;
   20982: out<=1;
   20983: out<=0;
   20984: out<=1;
   20985: out<=0;
   20986: out<=1;
   20987: out<=0;
   20988: out<=1;
   20989: out<=1;
   20990: out<=0;
   20991: out<=0;
   20992: out<=0;
   20993: out<=0;
   20994: out<=0;
   20995: out<=0;
   20996: out<=0;
   20997: out<=1;
   20998: out<=1;
   20999: out<=0;
   21000: out<=1;
   21001: out<=0;
   21002: out<=1;
   21003: out<=0;
   21004: out<=1;
   21005: out<=1;
   21006: out<=0;
   21007: out<=0;
   21008: out<=0;
   21009: out<=1;
   21010: out<=1;
   21011: out<=0;
   21012: out<=1;
   21013: out<=1;
   21014: out<=1;
   21015: out<=1;
   21016: out<=0;
   21017: out<=0;
   21018: out<=1;
   21019: out<=1;
   21020: out<=1;
   21021: out<=0;
   21022: out<=1;
   21023: out<=0;
   21024: out<=0;
   21025: out<=1;
   21026: out<=0;
   21027: out<=1;
   21028: out<=1;
   21029: out<=1;
   21030: out<=0;
   21031: out<=0;
   21032: out<=1;
   21033: out<=1;
   21034: out<=1;
   21035: out<=1;
   21036: out<=0;
   21037: out<=1;
   21038: out<=1;
   21039: out<=0;
   21040: out<=0;
   21041: out<=0;
   21042: out<=1;
   21043: out<=1;
   21044: out<=0;
   21045: out<=1;
   21046: out<=0;
   21047: out<=1;
   21048: out<=0;
   21049: out<=1;
   21050: out<=1;
   21051: out<=0;
   21052: out<=0;
   21053: out<=0;
   21054: out<=0;
   21055: out<=0;
   21056: out<=1;
   21057: out<=1;
   21058: out<=1;
   21059: out<=1;
   21060: out<=1;
   21061: out<=0;
   21062: out<=0;
   21063: out<=1;
   21064: out<=0;
   21065: out<=1;
   21066: out<=0;
   21067: out<=1;
   21068: out<=0;
   21069: out<=0;
   21070: out<=1;
   21071: out<=1;
   21072: out<=0;
   21073: out<=1;
   21074: out<=1;
   21075: out<=0;
   21076: out<=1;
   21077: out<=1;
   21078: out<=1;
   21079: out<=1;
   21080: out<=0;
   21081: out<=0;
   21082: out<=1;
   21083: out<=1;
   21084: out<=1;
   21085: out<=0;
   21086: out<=1;
   21087: out<=0;
   21088: out<=0;
   21089: out<=1;
   21090: out<=0;
   21091: out<=1;
   21092: out<=1;
   21093: out<=1;
   21094: out<=0;
   21095: out<=0;
   21096: out<=1;
   21097: out<=1;
   21098: out<=1;
   21099: out<=1;
   21100: out<=0;
   21101: out<=1;
   21102: out<=1;
   21103: out<=0;
   21104: out<=1;
   21105: out<=1;
   21106: out<=0;
   21107: out<=0;
   21108: out<=1;
   21109: out<=0;
   21110: out<=1;
   21111: out<=0;
   21112: out<=1;
   21113: out<=0;
   21114: out<=0;
   21115: out<=1;
   21116: out<=1;
   21117: out<=1;
   21118: out<=1;
   21119: out<=1;
   21120: out<=1;
   21121: out<=1;
   21122: out<=1;
   21123: out<=1;
   21124: out<=1;
   21125: out<=0;
   21126: out<=0;
   21127: out<=1;
   21128: out<=0;
   21129: out<=1;
   21130: out<=0;
   21131: out<=1;
   21132: out<=0;
   21133: out<=0;
   21134: out<=1;
   21135: out<=1;
   21136: out<=0;
   21137: out<=1;
   21138: out<=1;
   21139: out<=0;
   21140: out<=1;
   21141: out<=1;
   21142: out<=1;
   21143: out<=1;
   21144: out<=0;
   21145: out<=0;
   21146: out<=1;
   21147: out<=1;
   21148: out<=1;
   21149: out<=0;
   21150: out<=1;
   21151: out<=0;
   21152: out<=1;
   21153: out<=0;
   21154: out<=1;
   21155: out<=0;
   21156: out<=0;
   21157: out<=0;
   21158: out<=1;
   21159: out<=1;
   21160: out<=0;
   21161: out<=0;
   21162: out<=0;
   21163: out<=0;
   21164: out<=1;
   21165: out<=0;
   21166: out<=0;
   21167: out<=1;
   21168: out<=0;
   21169: out<=0;
   21170: out<=1;
   21171: out<=1;
   21172: out<=0;
   21173: out<=1;
   21174: out<=0;
   21175: out<=1;
   21176: out<=0;
   21177: out<=1;
   21178: out<=1;
   21179: out<=0;
   21180: out<=0;
   21181: out<=0;
   21182: out<=0;
   21183: out<=0;
   21184: out<=0;
   21185: out<=0;
   21186: out<=0;
   21187: out<=0;
   21188: out<=0;
   21189: out<=1;
   21190: out<=1;
   21191: out<=0;
   21192: out<=1;
   21193: out<=0;
   21194: out<=1;
   21195: out<=0;
   21196: out<=1;
   21197: out<=1;
   21198: out<=0;
   21199: out<=0;
   21200: out<=0;
   21201: out<=1;
   21202: out<=1;
   21203: out<=0;
   21204: out<=1;
   21205: out<=1;
   21206: out<=1;
   21207: out<=1;
   21208: out<=0;
   21209: out<=0;
   21210: out<=1;
   21211: out<=1;
   21212: out<=1;
   21213: out<=0;
   21214: out<=1;
   21215: out<=0;
   21216: out<=1;
   21217: out<=0;
   21218: out<=1;
   21219: out<=0;
   21220: out<=0;
   21221: out<=0;
   21222: out<=1;
   21223: out<=1;
   21224: out<=0;
   21225: out<=0;
   21226: out<=0;
   21227: out<=0;
   21228: out<=1;
   21229: out<=0;
   21230: out<=0;
   21231: out<=1;
   21232: out<=1;
   21233: out<=1;
   21234: out<=0;
   21235: out<=0;
   21236: out<=1;
   21237: out<=0;
   21238: out<=1;
   21239: out<=0;
   21240: out<=1;
   21241: out<=0;
   21242: out<=0;
   21243: out<=1;
   21244: out<=1;
   21245: out<=1;
   21246: out<=1;
   21247: out<=1;
   21248: out<=0;
   21249: out<=1;
   21250: out<=1;
   21251: out<=0;
   21252: out<=1;
   21253: out<=1;
   21254: out<=1;
   21255: out<=1;
   21256: out<=0;
   21257: out<=0;
   21258: out<=1;
   21259: out<=1;
   21260: out<=1;
   21261: out<=0;
   21262: out<=1;
   21263: out<=0;
   21264: out<=1;
   21265: out<=1;
   21266: out<=1;
   21267: out<=1;
   21268: out<=1;
   21269: out<=0;
   21270: out<=0;
   21271: out<=1;
   21272: out<=0;
   21273: out<=1;
   21274: out<=0;
   21275: out<=1;
   21276: out<=0;
   21277: out<=0;
   21278: out<=1;
   21279: out<=1;
   21280: out<=1;
   21281: out<=1;
   21282: out<=0;
   21283: out<=0;
   21284: out<=1;
   21285: out<=0;
   21286: out<=1;
   21287: out<=0;
   21288: out<=1;
   21289: out<=0;
   21290: out<=0;
   21291: out<=1;
   21292: out<=1;
   21293: out<=1;
   21294: out<=1;
   21295: out<=1;
   21296: out<=0;
   21297: out<=1;
   21298: out<=0;
   21299: out<=1;
   21300: out<=1;
   21301: out<=1;
   21302: out<=0;
   21303: out<=0;
   21304: out<=1;
   21305: out<=1;
   21306: out<=1;
   21307: out<=1;
   21308: out<=0;
   21309: out<=1;
   21310: out<=1;
   21311: out<=0;
   21312: out<=0;
   21313: out<=1;
   21314: out<=1;
   21315: out<=0;
   21316: out<=1;
   21317: out<=1;
   21318: out<=1;
   21319: out<=1;
   21320: out<=0;
   21321: out<=0;
   21322: out<=1;
   21323: out<=1;
   21324: out<=1;
   21325: out<=0;
   21326: out<=1;
   21327: out<=0;
   21328: out<=0;
   21329: out<=0;
   21330: out<=0;
   21331: out<=0;
   21332: out<=0;
   21333: out<=1;
   21334: out<=1;
   21335: out<=0;
   21336: out<=1;
   21337: out<=0;
   21338: out<=1;
   21339: out<=0;
   21340: out<=1;
   21341: out<=1;
   21342: out<=0;
   21343: out<=0;
   21344: out<=0;
   21345: out<=0;
   21346: out<=1;
   21347: out<=1;
   21348: out<=0;
   21349: out<=1;
   21350: out<=0;
   21351: out<=1;
   21352: out<=0;
   21353: out<=1;
   21354: out<=1;
   21355: out<=0;
   21356: out<=0;
   21357: out<=0;
   21358: out<=0;
   21359: out<=0;
   21360: out<=0;
   21361: out<=1;
   21362: out<=0;
   21363: out<=1;
   21364: out<=1;
   21365: out<=1;
   21366: out<=0;
   21367: out<=0;
   21368: out<=1;
   21369: out<=1;
   21370: out<=1;
   21371: out<=1;
   21372: out<=0;
   21373: out<=1;
   21374: out<=1;
   21375: out<=0;
   21376: out<=0;
   21377: out<=1;
   21378: out<=1;
   21379: out<=0;
   21380: out<=1;
   21381: out<=1;
   21382: out<=1;
   21383: out<=1;
   21384: out<=0;
   21385: out<=0;
   21386: out<=1;
   21387: out<=1;
   21388: out<=1;
   21389: out<=0;
   21390: out<=1;
   21391: out<=0;
   21392: out<=0;
   21393: out<=0;
   21394: out<=0;
   21395: out<=0;
   21396: out<=0;
   21397: out<=1;
   21398: out<=1;
   21399: out<=0;
   21400: out<=1;
   21401: out<=0;
   21402: out<=1;
   21403: out<=0;
   21404: out<=1;
   21405: out<=1;
   21406: out<=0;
   21407: out<=0;
   21408: out<=1;
   21409: out<=1;
   21410: out<=0;
   21411: out<=0;
   21412: out<=1;
   21413: out<=0;
   21414: out<=1;
   21415: out<=0;
   21416: out<=1;
   21417: out<=0;
   21418: out<=0;
   21419: out<=1;
   21420: out<=1;
   21421: out<=1;
   21422: out<=1;
   21423: out<=1;
   21424: out<=1;
   21425: out<=0;
   21426: out<=1;
   21427: out<=0;
   21428: out<=0;
   21429: out<=0;
   21430: out<=1;
   21431: out<=1;
   21432: out<=0;
   21433: out<=0;
   21434: out<=0;
   21435: out<=0;
   21436: out<=1;
   21437: out<=0;
   21438: out<=0;
   21439: out<=1;
   21440: out<=0;
   21441: out<=1;
   21442: out<=1;
   21443: out<=0;
   21444: out<=1;
   21445: out<=1;
   21446: out<=1;
   21447: out<=1;
   21448: out<=0;
   21449: out<=0;
   21450: out<=1;
   21451: out<=1;
   21452: out<=1;
   21453: out<=0;
   21454: out<=1;
   21455: out<=0;
   21456: out<=1;
   21457: out<=1;
   21458: out<=1;
   21459: out<=1;
   21460: out<=1;
   21461: out<=0;
   21462: out<=0;
   21463: out<=1;
   21464: out<=0;
   21465: out<=1;
   21466: out<=0;
   21467: out<=1;
   21468: out<=0;
   21469: out<=0;
   21470: out<=1;
   21471: out<=1;
   21472: out<=0;
   21473: out<=0;
   21474: out<=1;
   21475: out<=1;
   21476: out<=0;
   21477: out<=1;
   21478: out<=0;
   21479: out<=1;
   21480: out<=0;
   21481: out<=1;
   21482: out<=1;
   21483: out<=0;
   21484: out<=0;
   21485: out<=0;
   21486: out<=0;
   21487: out<=0;
   21488: out<=1;
   21489: out<=0;
   21490: out<=1;
   21491: out<=0;
   21492: out<=0;
   21493: out<=0;
   21494: out<=1;
   21495: out<=1;
   21496: out<=0;
   21497: out<=0;
   21498: out<=0;
   21499: out<=0;
   21500: out<=1;
   21501: out<=0;
   21502: out<=0;
   21503: out<=1;
   21504: out<=1;
   21505: out<=1;
   21506: out<=0;
   21507: out<=0;
   21508: out<=0;
   21509: out<=1;
   21510: out<=0;
   21511: out<=1;
   21512: out<=0;
   21513: out<=1;
   21514: out<=1;
   21515: out<=0;
   21516: out<=1;
   21517: out<=1;
   21518: out<=1;
   21519: out<=1;
   21520: out<=0;
   21521: out<=1;
   21522: out<=0;
   21523: out<=1;
   21524: out<=0;
   21525: out<=0;
   21526: out<=1;
   21527: out<=1;
   21528: out<=0;
   21529: out<=0;
   21530: out<=0;
   21531: out<=0;
   21532: out<=0;
   21533: out<=1;
   21534: out<=1;
   21535: out<=0;
   21536: out<=1;
   21537: out<=0;
   21538: out<=0;
   21539: out<=1;
   21540: out<=1;
   21541: out<=1;
   21542: out<=1;
   21543: out<=1;
   21544: out<=0;
   21545: out<=0;
   21546: out<=1;
   21547: out<=1;
   21548: out<=0;
   21549: out<=1;
   21550: out<=0;
   21551: out<=1;
   21552: out<=0;
   21553: out<=0;
   21554: out<=0;
   21555: out<=0;
   21556: out<=1;
   21557: out<=0;
   21558: out<=0;
   21559: out<=1;
   21560: out<=0;
   21561: out<=1;
   21562: out<=0;
   21563: out<=1;
   21564: out<=1;
   21565: out<=1;
   21566: out<=0;
   21567: out<=0;
   21568: out<=0;
   21569: out<=0;
   21570: out<=1;
   21571: out<=1;
   21572: out<=1;
   21573: out<=0;
   21574: out<=1;
   21575: out<=0;
   21576: out<=1;
   21577: out<=0;
   21578: out<=0;
   21579: out<=1;
   21580: out<=0;
   21581: out<=0;
   21582: out<=0;
   21583: out<=0;
   21584: out<=0;
   21585: out<=1;
   21586: out<=0;
   21587: out<=1;
   21588: out<=0;
   21589: out<=0;
   21590: out<=1;
   21591: out<=1;
   21592: out<=0;
   21593: out<=0;
   21594: out<=0;
   21595: out<=0;
   21596: out<=0;
   21597: out<=1;
   21598: out<=1;
   21599: out<=0;
   21600: out<=1;
   21601: out<=0;
   21602: out<=0;
   21603: out<=1;
   21604: out<=1;
   21605: out<=1;
   21606: out<=1;
   21607: out<=1;
   21608: out<=0;
   21609: out<=0;
   21610: out<=1;
   21611: out<=1;
   21612: out<=0;
   21613: out<=1;
   21614: out<=0;
   21615: out<=1;
   21616: out<=1;
   21617: out<=1;
   21618: out<=1;
   21619: out<=1;
   21620: out<=0;
   21621: out<=1;
   21622: out<=1;
   21623: out<=0;
   21624: out<=1;
   21625: out<=0;
   21626: out<=1;
   21627: out<=0;
   21628: out<=0;
   21629: out<=0;
   21630: out<=1;
   21631: out<=1;
   21632: out<=1;
   21633: out<=1;
   21634: out<=0;
   21635: out<=0;
   21636: out<=0;
   21637: out<=1;
   21638: out<=0;
   21639: out<=1;
   21640: out<=0;
   21641: out<=1;
   21642: out<=1;
   21643: out<=0;
   21644: out<=1;
   21645: out<=1;
   21646: out<=1;
   21647: out<=1;
   21648: out<=1;
   21649: out<=0;
   21650: out<=1;
   21651: out<=0;
   21652: out<=1;
   21653: out<=1;
   21654: out<=0;
   21655: out<=0;
   21656: out<=1;
   21657: out<=1;
   21658: out<=1;
   21659: out<=1;
   21660: out<=1;
   21661: out<=0;
   21662: out<=0;
   21663: out<=1;
   21664: out<=1;
   21665: out<=0;
   21666: out<=0;
   21667: out<=1;
   21668: out<=1;
   21669: out<=1;
   21670: out<=1;
   21671: out<=1;
   21672: out<=0;
   21673: out<=0;
   21674: out<=1;
   21675: out<=1;
   21676: out<=0;
   21677: out<=1;
   21678: out<=0;
   21679: out<=1;
   21680: out<=1;
   21681: out<=1;
   21682: out<=1;
   21683: out<=1;
   21684: out<=0;
   21685: out<=1;
   21686: out<=1;
   21687: out<=0;
   21688: out<=1;
   21689: out<=0;
   21690: out<=1;
   21691: out<=0;
   21692: out<=0;
   21693: out<=0;
   21694: out<=1;
   21695: out<=1;
   21696: out<=0;
   21697: out<=0;
   21698: out<=1;
   21699: out<=1;
   21700: out<=1;
   21701: out<=0;
   21702: out<=1;
   21703: out<=0;
   21704: out<=1;
   21705: out<=0;
   21706: out<=0;
   21707: out<=1;
   21708: out<=0;
   21709: out<=0;
   21710: out<=0;
   21711: out<=0;
   21712: out<=1;
   21713: out<=0;
   21714: out<=1;
   21715: out<=0;
   21716: out<=1;
   21717: out<=1;
   21718: out<=0;
   21719: out<=0;
   21720: out<=1;
   21721: out<=1;
   21722: out<=1;
   21723: out<=1;
   21724: out<=1;
   21725: out<=0;
   21726: out<=0;
   21727: out<=1;
   21728: out<=1;
   21729: out<=0;
   21730: out<=0;
   21731: out<=1;
   21732: out<=1;
   21733: out<=1;
   21734: out<=1;
   21735: out<=1;
   21736: out<=0;
   21737: out<=0;
   21738: out<=1;
   21739: out<=1;
   21740: out<=0;
   21741: out<=1;
   21742: out<=0;
   21743: out<=1;
   21744: out<=0;
   21745: out<=0;
   21746: out<=0;
   21747: out<=0;
   21748: out<=1;
   21749: out<=0;
   21750: out<=0;
   21751: out<=1;
   21752: out<=0;
   21753: out<=1;
   21754: out<=0;
   21755: out<=1;
   21756: out<=1;
   21757: out<=1;
   21758: out<=0;
   21759: out<=0;
   21760: out<=0;
   21761: out<=1;
   21762: out<=0;
   21763: out<=1;
   21764: out<=0;
   21765: out<=0;
   21766: out<=1;
   21767: out<=1;
   21768: out<=0;
   21769: out<=0;
   21770: out<=0;
   21771: out<=0;
   21772: out<=0;
   21773: out<=1;
   21774: out<=1;
   21775: out<=0;
   21776: out<=0;
   21777: out<=0;
   21778: out<=1;
   21779: out<=1;
   21780: out<=1;
   21781: out<=0;
   21782: out<=1;
   21783: out<=0;
   21784: out<=1;
   21785: out<=0;
   21786: out<=0;
   21787: out<=1;
   21788: out<=0;
   21789: out<=0;
   21790: out<=0;
   21791: out<=0;
   21792: out<=1;
   21793: out<=1;
   21794: out<=1;
   21795: out<=1;
   21796: out<=0;
   21797: out<=1;
   21798: out<=1;
   21799: out<=0;
   21800: out<=1;
   21801: out<=0;
   21802: out<=1;
   21803: out<=0;
   21804: out<=0;
   21805: out<=0;
   21806: out<=1;
   21807: out<=1;
   21808: out<=1;
   21809: out<=0;
   21810: out<=0;
   21811: out<=1;
   21812: out<=1;
   21813: out<=1;
   21814: out<=1;
   21815: out<=1;
   21816: out<=0;
   21817: out<=0;
   21818: out<=1;
   21819: out<=1;
   21820: out<=0;
   21821: out<=1;
   21822: out<=0;
   21823: out<=1;
   21824: out<=0;
   21825: out<=1;
   21826: out<=0;
   21827: out<=1;
   21828: out<=0;
   21829: out<=0;
   21830: out<=1;
   21831: out<=1;
   21832: out<=0;
   21833: out<=0;
   21834: out<=0;
   21835: out<=0;
   21836: out<=0;
   21837: out<=1;
   21838: out<=1;
   21839: out<=0;
   21840: out<=1;
   21841: out<=1;
   21842: out<=0;
   21843: out<=0;
   21844: out<=0;
   21845: out<=1;
   21846: out<=0;
   21847: out<=1;
   21848: out<=0;
   21849: out<=1;
   21850: out<=1;
   21851: out<=0;
   21852: out<=1;
   21853: out<=1;
   21854: out<=1;
   21855: out<=1;
   21856: out<=0;
   21857: out<=0;
   21858: out<=0;
   21859: out<=0;
   21860: out<=1;
   21861: out<=0;
   21862: out<=0;
   21863: out<=1;
   21864: out<=0;
   21865: out<=1;
   21866: out<=0;
   21867: out<=1;
   21868: out<=1;
   21869: out<=1;
   21870: out<=0;
   21871: out<=0;
   21872: out<=1;
   21873: out<=0;
   21874: out<=0;
   21875: out<=1;
   21876: out<=1;
   21877: out<=1;
   21878: out<=1;
   21879: out<=1;
   21880: out<=0;
   21881: out<=0;
   21882: out<=1;
   21883: out<=1;
   21884: out<=0;
   21885: out<=1;
   21886: out<=0;
   21887: out<=1;
   21888: out<=1;
   21889: out<=0;
   21890: out<=1;
   21891: out<=0;
   21892: out<=1;
   21893: out<=1;
   21894: out<=0;
   21895: out<=0;
   21896: out<=1;
   21897: out<=1;
   21898: out<=1;
   21899: out<=1;
   21900: out<=1;
   21901: out<=0;
   21902: out<=0;
   21903: out<=1;
   21904: out<=0;
   21905: out<=0;
   21906: out<=1;
   21907: out<=1;
   21908: out<=1;
   21909: out<=0;
   21910: out<=1;
   21911: out<=0;
   21912: out<=1;
   21913: out<=0;
   21914: out<=0;
   21915: out<=1;
   21916: out<=0;
   21917: out<=0;
   21918: out<=0;
   21919: out<=0;
   21920: out<=0;
   21921: out<=0;
   21922: out<=0;
   21923: out<=0;
   21924: out<=1;
   21925: out<=0;
   21926: out<=0;
   21927: out<=1;
   21928: out<=0;
   21929: out<=1;
   21930: out<=0;
   21931: out<=1;
   21932: out<=1;
   21933: out<=1;
   21934: out<=0;
   21935: out<=0;
   21936: out<=1;
   21937: out<=0;
   21938: out<=0;
   21939: out<=1;
   21940: out<=1;
   21941: out<=1;
   21942: out<=1;
   21943: out<=1;
   21944: out<=0;
   21945: out<=0;
   21946: out<=1;
   21947: out<=1;
   21948: out<=0;
   21949: out<=1;
   21950: out<=0;
   21951: out<=1;
   21952: out<=1;
   21953: out<=0;
   21954: out<=1;
   21955: out<=0;
   21956: out<=1;
   21957: out<=1;
   21958: out<=0;
   21959: out<=0;
   21960: out<=1;
   21961: out<=1;
   21962: out<=1;
   21963: out<=1;
   21964: out<=1;
   21965: out<=0;
   21966: out<=0;
   21967: out<=1;
   21968: out<=1;
   21969: out<=1;
   21970: out<=0;
   21971: out<=0;
   21972: out<=0;
   21973: out<=1;
   21974: out<=0;
   21975: out<=1;
   21976: out<=0;
   21977: out<=1;
   21978: out<=1;
   21979: out<=0;
   21980: out<=1;
   21981: out<=1;
   21982: out<=1;
   21983: out<=1;
   21984: out<=1;
   21985: out<=1;
   21986: out<=1;
   21987: out<=1;
   21988: out<=0;
   21989: out<=1;
   21990: out<=1;
   21991: out<=0;
   21992: out<=1;
   21993: out<=0;
   21994: out<=1;
   21995: out<=0;
   21996: out<=0;
   21997: out<=0;
   21998: out<=1;
   21999: out<=1;
   22000: out<=1;
   22001: out<=0;
   22002: out<=0;
   22003: out<=1;
   22004: out<=1;
   22005: out<=1;
   22006: out<=1;
   22007: out<=1;
   22008: out<=0;
   22009: out<=0;
   22010: out<=1;
   22011: out<=1;
   22012: out<=0;
   22013: out<=1;
   22014: out<=0;
   22015: out<=1;
   22016: out<=1;
   22017: out<=0;
   22018: out<=0;
   22019: out<=1;
   22020: out<=1;
   22021: out<=1;
   22022: out<=1;
   22023: out<=1;
   22024: out<=0;
   22025: out<=0;
   22026: out<=1;
   22027: out<=1;
   22028: out<=0;
   22029: out<=1;
   22030: out<=0;
   22031: out<=1;
   22032: out<=1;
   22033: out<=1;
   22034: out<=1;
   22035: out<=1;
   22036: out<=0;
   22037: out<=1;
   22038: out<=1;
   22039: out<=0;
   22040: out<=1;
   22041: out<=0;
   22042: out<=1;
   22043: out<=0;
   22044: out<=0;
   22045: out<=0;
   22046: out<=1;
   22047: out<=1;
   22048: out<=1;
   22049: out<=1;
   22050: out<=0;
   22051: out<=0;
   22052: out<=0;
   22053: out<=1;
   22054: out<=0;
   22055: out<=1;
   22056: out<=0;
   22057: out<=1;
   22058: out<=1;
   22059: out<=0;
   22060: out<=1;
   22061: out<=1;
   22062: out<=1;
   22063: out<=1;
   22064: out<=1;
   22065: out<=0;
   22066: out<=1;
   22067: out<=0;
   22068: out<=1;
   22069: out<=1;
   22070: out<=0;
   22071: out<=0;
   22072: out<=1;
   22073: out<=1;
   22074: out<=1;
   22075: out<=1;
   22076: out<=1;
   22077: out<=0;
   22078: out<=0;
   22079: out<=1;
   22080: out<=1;
   22081: out<=0;
   22082: out<=0;
   22083: out<=1;
   22084: out<=1;
   22085: out<=1;
   22086: out<=1;
   22087: out<=1;
   22088: out<=0;
   22089: out<=0;
   22090: out<=1;
   22091: out<=1;
   22092: out<=0;
   22093: out<=1;
   22094: out<=0;
   22095: out<=1;
   22096: out<=0;
   22097: out<=0;
   22098: out<=0;
   22099: out<=0;
   22100: out<=1;
   22101: out<=0;
   22102: out<=0;
   22103: out<=1;
   22104: out<=0;
   22105: out<=1;
   22106: out<=0;
   22107: out<=1;
   22108: out<=1;
   22109: out<=1;
   22110: out<=0;
   22111: out<=0;
   22112: out<=0;
   22113: out<=0;
   22114: out<=1;
   22115: out<=1;
   22116: out<=1;
   22117: out<=0;
   22118: out<=1;
   22119: out<=0;
   22120: out<=1;
   22121: out<=0;
   22122: out<=0;
   22123: out<=1;
   22124: out<=0;
   22125: out<=0;
   22126: out<=0;
   22127: out<=0;
   22128: out<=1;
   22129: out<=0;
   22130: out<=1;
   22131: out<=0;
   22132: out<=1;
   22133: out<=1;
   22134: out<=0;
   22135: out<=0;
   22136: out<=1;
   22137: out<=1;
   22138: out<=1;
   22139: out<=1;
   22140: out<=1;
   22141: out<=0;
   22142: out<=0;
   22143: out<=1;
   22144: out<=1;
   22145: out<=0;
   22146: out<=0;
   22147: out<=1;
   22148: out<=1;
   22149: out<=1;
   22150: out<=1;
   22151: out<=1;
   22152: out<=0;
   22153: out<=0;
   22154: out<=1;
   22155: out<=1;
   22156: out<=0;
   22157: out<=1;
   22158: out<=0;
   22159: out<=1;
   22160: out<=0;
   22161: out<=0;
   22162: out<=0;
   22163: out<=0;
   22164: out<=1;
   22165: out<=0;
   22166: out<=0;
   22167: out<=1;
   22168: out<=0;
   22169: out<=1;
   22170: out<=0;
   22171: out<=1;
   22172: out<=1;
   22173: out<=1;
   22174: out<=0;
   22175: out<=0;
   22176: out<=1;
   22177: out<=1;
   22178: out<=0;
   22179: out<=0;
   22180: out<=0;
   22181: out<=1;
   22182: out<=0;
   22183: out<=1;
   22184: out<=0;
   22185: out<=1;
   22186: out<=1;
   22187: out<=0;
   22188: out<=1;
   22189: out<=1;
   22190: out<=1;
   22191: out<=1;
   22192: out<=0;
   22193: out<=1;
   22194: out<=0;
   22195: out<=1;
   22196: out<=0;
   22197: out<=0;
   22198: out<=1;
   22199: out<=1;
   22200: out<=0;
   22201: out<=0;
   22202: out<=0;
   22203: out<=0;
   22204: out<=0;
   22205: out<=1;
   22206: out<=1;
   22207: out<=0;
   22208: out<=1;
   22209: out<=0;
   22210: out<=0;
   22211: out<=1;
   22212: out<=1;
   22213: out<=1;
   22214: out<=1;
   22215: out<=1;
   22216: out<=0;
   22217: out<=0;
   22218: out<=1;
   22219: out<=1;
   22220: out<=0;
   22221: out<=1;
   22222: out<=0;
   22223: out<=1;
   22224: out<=1;
   22225: out<=1;
   22226: out<=1;
   22227: out<=1;
   22228: out<=0;
   22229: out<=1;
   22230: out<=1;
   22231: out<=0;
   22232: out<=1;
   22233: out<=0;
   22234: out<=1;
   22235: out<=0;
   22236: out<=0;
   22237: out<=0;
   22238: out<=1;
   22239: out<=1;
   22240: out<=0;
   22241: out<=0;
   22242: out<=1;
   22243: out<=1;
   22244: out<=1;
   22245: out<=0;
   22246: out<=1;
   22247: out<=0;
   22248: out<=1;
   22249: out<=0;
   22250: out<=0;
   22251: out<=1;
   22252: out<=0;
   22253: out<=0;
   22254: out<=0;
   22255: out<=0;
   22256: out<=0;
   22257: out<=1;
   22258: out<=0;
   22259: out<=1;
   22260: out<=0;
   22261: out<=0;
   22262: out<=1;
   22263: out<=1;
   22264: out<=0;
   22265: out<=0;
   22266: out<=0;
   22267: out<=0;
   22268: out<=0;
   22269: out<=1;
   22270: out<=1;
   22271: out<=0;
   22272: out<=0;
   22273: out<=0;
   22274: out<=0;
   22275: out<=0;
   22276: out<=1;
   22277: out<=0;
   22278: out<=0;
   22279: out<=1;
   22280: out<=0;
   22281: out<=1;
   22282: out<=0;
   22283: out<=1;
   22284: out<=1;
   22285: out<=1;
   22286: out<=0;
   22287: out<=0;
   22288: out<=1;
   22289: out<=0;
   22290: out<=0;
   22291: out<=1;
   22292: out<=1;
   22293: out<=1;
   22294: out<=1;
   22295: out<=1;
   22296: out<=0;
   22297: out<=0;
   22298: out<=1;
   22299: out<=1;
   22300: out<=0;
   22301: out<=1;
   22302: out<=0;
   22303: out<=1;
   22304: out<=1;
   22305: out<=0;
   22306: out<=1;
   22307: out<=0;
   22308: out<=1;
   22309: out<=1;
   22310: out<=0;
   22311: out<=0;
   22312: out<=1;
   22313: out<=1;
   22314: out<=1;
   22315: out<=1;
   22316: out<=1;
   22317: out<=0;
   22318: out<=0;
   22319: out<=1;
   22320: out<=0;
   22321: out<=0;
   22322: out<=1;
   22323: out<=1;
   22324: out<=1;
   22325: out<=0;
   22326: out<=1;
   22327: out<=0;
   22328: out<=1;
   22329: out<=0;
   22330: out<=0;
   22331: out<=1;
   22332: out<=0;
   22333: out<=0;
   22334: out<=0;
   22335: out<=0;
   22336: out<=1;
   22337: out<=1;
   22338: out<=1;
   22339: out<=1;
   22340: out<=0;
   22341: out<=1;
   22342: out<=1;
   22343: out<=0;
   22344: out<=1;
   22345: out<=0;
   22346: out<=1;
   22347: out<=0;
   22348: out<=0;
   22349: out<=0;
   22350: out<=1;
   22351: out<=1;
   22352: out<=1;
   22353: out<=0;
   22354: out<=0;
   22355: out<=1;
   22356: out<=1;
   22357: out<=1;
   22358: out<=1;
   22359: out<=1;
   22360: out<=0;
   22361: out<=0;
   22362: out<=1;
   22363: out<=1;
   22364: out<=0;
   22365: out<=1;
   22366: out<=0;
   22367: out<=1;
   22368: out<=1;
   22369: out<=0;
   22370: out<=1;
   22371: out<=0;
   22372: out<=1;
   22373: out<=1;
   22374: out<=0;
   22375: out<=0;
   22376: out<=1;
   22377: out<=1;
   22378: out<=1;
   22379: out<=1;
   22380: out<=1;
   22381: out<=0;
   22382: out<=0;
   22383: out<=1;
   22384: out<=1;
   22385: out<=1;
   22386: out<=0;
   22387: out<=0;
   22388: out<=0;
   22389: out<=1;
   22390: out<=0;
   22391: out<=1;
   22392: out<=0;
   22393: out<=1;
   22394: out<=1;
   22395: out<=0;
   22396: out<=1;
   22397: out<=1;
   22398: out<=1;
   22399: out<=1;
   22400: out<=1;
   22401: out<=1;
   22402: out<=1;
   22403: out<=1;
   22404: out<=0;
   22405: out<=1;
   22406: out<=1;
   22407: out<=0;
   22408: out<=1;
   22409: out<=0;
   22410: out<=1;
   22411: out<=0;
   22412: out<=0;
   22413: out<=0;
   22414: out<=1;
   22415: out<=1;
   22416: out<=1;
   22417: out<=0;
   22418: out<=0;
   22419: out<=1;
   22420: out<=1;
   22421: out<=1;
   22422: out<=1;
   22423: out<=1;
   22424: out<=0;
   22425: out<=0;
   22426: out<=1;
   22427: out<=1;
   22428: out<=0;
   22429: out<=1;
   22430: out<=0;
   22431: out<=1;
   22432: out<=0;
   22433: out<=1;
   22434: out<=0;
   22435: out<=1;
   22436: out<=0;
   22437: out<=0;
   22438: out<=1;
   22439: out<=1;
   22440: out<=0;
   22441: out<=0;
   22442: out<=0;
   22443: out<=0;
   22444: out<=0;
   22445: out<=1;
   22446: out<=1;
   22447: out<=0;
   22448: out<=0;
   22449: out<=0;
   22450: out<=1;
   22451: out<=1;
   22452: out<=1;
   22453: out<=0;
   22454: out<=1;
   22455: out<=0;
   22456: out<=1;
   22457: out<=0;
   22458: out<=0;
   22459: out<=1;
   22460: out<=0;
   22461: out<=0;
   22462: out<=0;
   22463: out<=0;
   22464: out<=0;
   22465: out<=0;
   22466: out<=0;
   22467: out<=0;
   22468: out<=1;
   22469: out<=0;
   22470: out<=0;
   22471: out<=1;
   22472: out<=0;
   22473: out<=1;
   22474: out<=0;
   22475: out<=1;
   22476: out<=1;
   22477: out<=1;
   22478: out<=0;
   22479: out<=0;
   22480: out<=1;
   22481: out<=0;
   22482: out<=0;
   22483: out<=1;
   22484: out<=1;
   22485: out<=1;
   22486: out<=1;
   22487: out<=1;
   22488: out<=0;
   22489: out<=0;
   22490: out<=1;
   22491: out<=1;
   22492: out<=0;
   22493: out<=1;
   22494: out<=0;
   22495: out<=1;
   22496: out<=0;
   22497: out<=1;
   22498: out<=0;
   22499: out<=1;
   22500: out<=0;
   22501: out<=0;
   22502: out<=1;
   22503: out<=1;
   22504: out<=0;
   22505: out<=0;
   22506: out<=0;
   22507: out<=0;
   22508: out<=0;
   22509: out<=1;
   22510: out<=1;
   22511: out<=0;
   22512: out<=1;
   22513: out<=1;
   22514: out<=0;
   22515: out<=0;
   22516: out<=0;
   22517: out<=1;
   22518: out<=0;
   22519: out<=1;
   22520: out<=0;
   22521: out<=1;
   22522: out<=1;
   22523: out<=0;
   22524: out<=1;
   22525: out<=1;
   22526: out<=1;
   22527: out<=1;
   22528: out<=0;
   22529: out<=0;
   22530: out<=0;
   22531: out<=0;
   22532: out<=1;
   22533: out<=0;
   22534: out<=0;
   22535: out<=1;
   22536: out<=1;
   22537: out<=0;
   22538: out<=1;
   22539: out<=0;
   22540: out<=0;
   22541: out<=0;
   22542: out<=1;
   22543: out<=1;
   22544: out<=1;
   22545: out<=0;
   22546: out<=0;
   22547: out<=1;
   22548: out<=1;
   22549: out<=1;
   22550: out<=1;
   22551: out<=1;
   22552: out<=1;
   22553: out<=1;
   22554: out<=0;
   22555: out<=0;
   22556: out<=1;
   22557: out<=0;
   22558: out<=1;
   22559: out<=0;
   22560: out<=0;
   22561: out<=1;
   22562: out<=0;
   22563: out<=1;
   22564: out<=0;
   22565: out<=0;
   22566: out<=1;
   22567: out<=1;
   22568: out<=1;
   22569: out<=1;
   22570: out<=1;
   22571: out<=1;
   22572: out<=1;
   22573: out<=0;
   22574: out<=0;
   22575: out<=1;
   22576: out<=1;
   22577: out<=1;
   22578: out<=0;
   22579: out<=0;
   22580: out<=0;
   22581: out<=1;
   22582: out<=0;
   22583: out<=1;
   22584: out<=1;
   22585: out<=0;
   22586: out<=0;
   22587: out<=1;
   22588: out<=0;
   22589: out<=0;
   22590: out<=0;
   22591: out<=0;
   22592: out<=1;
   22593: out<=1;
   22594: out<=1;
   22595: out<=1;
   22596: out<=0;
   22597: out<=1;
   22598: out<=1;
   22599: out<=0;
   22600: out<=0;
   22601: out<=1;
   22602: out<=0;
   22603: out<=1;
   22604: out<=1;
   22605: out<=1;
   22606: out<=0;
   22607: out<=0;
   22608: out<=1;
   22609: out<=0;
   22610: out<=0;
   22611: out<=1;
   22612: out<=1;
   22613: out<=1;
   22614: out<=1;
   22615: out<=1;
   22616: out<=1;
   22617: out<=1;
   22618: out<=0;
   22619: out<=0;
   22620: out<=1;
   22621: out<=0;
   22622: out<=1;
   22623: out<=0;
   22624: out<=0;
   22625: out<=1;
   22626: out<=0;
   22627: out<=1;
   22628: out<=0;
   22629: out<=0;
   22630: out<=1;
   22631: out<=1;
   22632: out<=1;
   22633: out<=1;
   22634: out<=1;
   22635: out<=1;
   22636: out<=1;
   22637: out<=0;
   22638: out<=0;
   22639: out<=1;
   22640: out<=0;
   22641: out<=0;
   22642: out<=1;
   22643: out<=1;
   22644: out<=1;
   22645: out<=0;
   22646: out<=1;
   22647: out<=0;
   22648: out<=0;
   22649: out<=1;
   22650: out<=1;
   22651: out<=0;
   22652: out<=1;
   22653: out<=1;
   22654: out<=1;
   22655: out<=1;
   22656: out<=1;
   22657: out<=1;
   22658: out<=1;
   22659: out<=1;
   22660: out<=0;
   22661: out<=1;
   22662: out<=1;
   22663: out<=0;
   22664: out<=0;
   22665: out<=1;
   22666: out<=0;
   22667: out<=1;
   22668: out<=1;
   22669: out<=1;
   22670: out<=0;
   22671: out<=0;
   22672: out<=1;
   22673: out<=0;
   22674: out<=0;
   22675: out<=1;
   22676: out<=1;
   22677: out<=1;
   22678: out<=1;
   22679: out<=1;
   22680: out<=1;
   22681: out<=1;
   22682: out<=0;
   22683: out<=0;
   22684: out<=1;
   22685: out<=0;
   22686: out<=1;
   22687: out<=0;
   22688: out<=1;
   22689: out<=0;
   22690: out<=1;
   22691: out<=0;
   22692: out<=1;
   22693: out<=1;
   22694: out<=0;
   22695: out<=0;
   22696: out<=0;
   22697: out<=0;
   22698: out<=0;
   22699: out<=0;
   22700: out<=0;
   22701: out<=1;
   22702: out<=1;
   22703: out<=0;
   22704: out<=1;
   22705: out<=1;
   22706: out<=0;
   22707: out<=0;
   22708: out<=0;
   22709: out<=1;
   22710: out<=0;
   22711: out<=1;
   22712: out<=1;
   22713: out<=0;
   22714: out<=0;
   22715: out<=1;
   22716: out<=0;
   22717: out<=0;
   22718: out<=0;
   22719: out<=0;
   22720: out<=0;
   22721: out<=0;
   22722: out<=0;
   22723: out<=0;
   22724: out<=1;
   22725: out<=0;
   22726: out<=0;
   22727: out<=1;
   22728: out<=1;
   22729: out<=0;
   22730: out<=1;
   22731: out<=0;
   22732: out<=0;
   22733: out<=0;
   22734: out<=1;
   22735: out<=1;
   22736: out<=1;
   22737: out<=0;
   22738: out<=0;
   22739: out<=1;
   22740: out<=1;
   22741: out<=1;
   22742: out<=1;
   22743: out<=1;
   22744: out<=1;
   22745: out<=1;
   22746: out<=0;
   22747: out<=0;
   22748: out<=1;
   22749: out<=0;
   22750: out<=1;
   22751: out<=0;
   22752: out<=1;
   22753: out<=0;
   22754: out<=1;
   22755: out<=0;
   22756: out<=1;
   22757: out<=1;
   22758: out<=0;
   22759: out<=0;
   22760: out<=0;
   22761: out<=0;
   22762: out<=0;
   22763: out<=0;
   22764: out<=0;
   22765: out<=1;
   22766: out<=1;
   22767: out<=0;
   22768: out<=0;
   22769: out<=0;
   22770: out<=1;
   22771: out<=1;
   22772: out<=1;
   22773: out<=0;
   22774: out<=1;
   22775: out<=0;
   22776: out<=0;
   22777: out<=1;
   22778: out<=1;
   22779: out<=0;
   22780: out<=1;
   22781: out<=1;
   22782: out<=1;
   22783: out<=1;
   22784: out<=1;
   22785: out<=0;
   22786: out<=0;
   22787: out<=1;
   22788: out<=1;
   22789: out<=1;
   22790: out<=1;
   22791: out<=1;
   22792: out<=1;
   22793: out<=1;
   22794: out<=0;
   22795: out<=0;
   22796: out<=1;
   22797: out<=0;
   22798: out<=1;
   22799: out<=0;
   22800: out<=1;
   22801: out<=1;
   22802: out<=1;
   22803: out<=1;
   22804: out<=0;
   22805: out<=1;
   22806: out<=1;
   22807: out<=0;
   22808: out<=0;
   22809: out<=1;
   22810: out<=0;
   22811: out<=1;
   22812: out<=1;
   22813: out<=1;
   22814: out<=0;
   22815: out<=0;
   22816: out<=0;
   22817: out<=0;
   22818: out<=1;
   22819: out<=1;
   22820: out<=1;
   22821: out<=0;
   22822: out<=1;
   22823: out<=0;
   22824: out<=0;
   22825: out<=1;
   22826: out<=1;
   22827: out<=0;
   22828: out<=1;
   22829: out<=1;
   22830: out<=1;
   22831: out<=1;
   22832: out<=0;
   22833: out<=1;
   22834: out<=0;
   22835: out<=1;
   22836: out<=0;
   22837: out<=0;
   22838: out<=1;
   22839: out<=1;
   22840: out<=1;
   22841: out<=1;
   22842: out<=1;
   22843: out<=1;
   22844: out<=1;
   22845: out<=0;
   22846: out<=0;
   22847: out<=1;
   22848: out<=1;
   22849: out<=0;
   22850: out<=0;
   22851: out<=1;
   22852: out<=1;
   22853: out<=1;
   22854: out<=1;
   22855: out<=1;
   22856: out<=1;
   22857: out<=1;
   22858: out<=0;
   22859: out<=0;
   22860: out<=1;
   22861: out<=0;
   22862: out<=1;
   22863: out<=0;
   22864: out<=0;
   22865: out<=0;
   22866: out<=0;
   22867: out<=0;
   22868: out<=1;
   22869: out<=0;
   22870: out<=0;
   22871: out<=1;
   22872: out<=1;
   22873: out<=0;
   22874: out<=1;
   22875: out<=0;
   22876: out<=0;
   22877: out<=0;
   22878: out<=1;
   22879: out<=1;
   22880: out<=1;
   22881: out<=1;
   22882: out<=0;
   22883: out<=0;
   22884: out<=0;
   22885: out<=1;
   22886: out<=0;
   22887: out<=1;
   22888: out<=1;
   22889: out<=0;
   22890: out<=0;
   22891: out<=1;
   22892: out<=0;
   22893: out<=0;
   22894: out<=0;
   22895: out<=0;
   22896: out<=0;
   22897: out<=1;
   22898: out<=0;
   22899: out<=1;
   22900: out<=0;
   22901: out<=0;
   22902: out<=1;
   22903: out<=1;
   22904: out<=1;
   22905: out<=1;
   22906: out<=1;
   22907: out<=1;
   22908: out<=1;
   22909: out<=0;
   22910: out<=0;
   22911: out<=1;
   22912: out<=1;
   22913: out<=0;
   22914: out<=0;
   22915: out<=1;
   22916: out<=1;
   22917: out<=1;
   22918: out<=1;
   22919: out<=1;
   22920: out<=1;
   22921: out<=1;
   22922: out<=0;
   22923: out<=0;
   22924: out<=1;
   22925: out<=0;
   22926: out<=1;
   22927: out<=0;
   22928: out<=0;
   22929: out<=0;
   22930: out<=0;
   22931: out<=0;
   22932: out<=1;
   22933: out<=0;
   22934: out<=0;
   22935: out<=1;
   22936: out<=1;
   22937: out<=0;
   22938: out<=1;
   22939: out<=0;
   22940: out<=0;
   22941: out<=0;
   22942: out<=1;
   22943: out<=1;
   22944: out<=0;
   22945: out<=0;
   22946: out<=1;
   22947: out<=1;
   22948: out<=1;
   22949: out<=0;
   22950: out<=1;
   22951: out<=0;
   22952: out<=0;
   22953: out<=1;
   22954: out<=1;
   22955: out<=0;
   22956: out<=1;
   22957: out<=1;
   22958: out<=1;
   22959: out<=1;
   22960: out<=1;
   22961: out<=0;
   22962: out<=1;
   22963: out<=0;
   22964: out<=1;
   22965: out<=1;
   22966: out<=0;
   22967: out<=0;
   22968: out<=0;
   22969: out<=0;
   22970: out<=0;
   22971: out<=0;
   22972: out<=0;
   22973: out<=1;
   22974: out<=1;
   22975: out<=0;
   22976: out<=1;
   22977: out<=0;
   22978: out<=0;
   22979: out<=1;
   22980: out<=1;
   22981: out<=1;
   22982: out<=1;
   22983: out<=1;
   22984: out<=1;
   22985: out<=1;
   22986: out<=0;
   22987: out<=0;
   22988: out<=1;
   22989: out<=0;
   22990: out<=1;
   22991: out<=0;
   22992: out<=1;
   22993: out<=1;
   22994: out<=1;
   22995: out<=1;
   22996: out<=0;
   22997: out<=1;
   22998: out<=1;
   22999: out<=0;
   23000: out<=0;
   23001: out<=1;
   23002: out<=0;
   23003: out<=1;
   23004: out<=1;
   23005: out<=1;
   23006: out<=0;
   23007: out<=0;
   23008: out<=1;
   23009: out<=1;
   23010: out<=0;
   23011: out<=0;
   23012: out<=0;
   23013: out<=1;
   23014: out<=0;
   23015: out<=1;
   23016: out<=1;
   23017: out<=0;
   23018: out<=0;
   23019: out<=1;
   23020: out<=0;
   23021: out<=0;
   23022: out<=0;
   23023: out<=0;
   23024: out<=1;
   23025: out<=0;
   23026: out<=1;
   23027: out<=0;
   23028: out<=1;
   23029: out<=1;
   23030: out<=0;
   23031: out<=0;
   23032: out<=0;
   23033: out<=0;
   23034: out<=0;
   23035: out<=0;
   23036: out<=0;
   23037: out<=1;
   23038: out<=1;
   23039: out<=0;
   23040: out<=1;
   23041: out<=0;
   23042: out<=1;
   23043: out<=0;
   23044: out<=1;
   23045: out<=1;
   23046: out<=0;
   23047: out<=0;
   23048: out<=0;
   23049: out<=0;
   23050: out<=0;
   23051: out<=0;
   23052: out<=0;
   23053: out<=1;
   23054: out<=1;
   23055: out<=0;
   23056: out<=1;
   23057: out<=1;
   23058: out<=0;
   23059: out<=0;
   23060: out<=0;
   23061: out<=1;
   23062: out<=0;
   23063: out<=1;
   23064: out<=1;
   23065: out<=0;
   23066: out<=0;
   23067: out<=1;
   23068: out<=0;
   23069: out<=0;
   23070: out<=0;
   23071: out<=0;
   23072: out<=1;
   23073: out<=1;
   23074: out<=1;
   23075: out<=1;
   23076: out<=0;
   23077: out<=1;
   23078: out<=1;
   23079: out<=0;
   23080: out<=0;
   23081: out<=1;
   23082: out<=0;
   23083: out<=1;
   23084: out<=1;
   23085: out<=1;
   23086: out<=0;
   23087: out<=0;
   23088: out<=1;
   23089: out<=0;
   23090: out<=0;
   23091: out<=1;
   23092: out<=1;
   23093: out<=1;
   23094: out<=1;
   23095: out<=1;
   23096: out<=1;
   23097: out<=1;
   23098: out<=0;
   23099: out<=0;
   23100: out<=1;
   23101: out<=0;
   23102: out<=1;
   23103: out<=0;
   23104: out<=1;
   23105: out<=0;
   23106: out<=1;
   23107: out<=0;
   23108: out<=1;
   23109: out<=1;
   23110: out<=0;
   23111: out<=0;
   23112: out<=0;
   23113: out<=0;
   23114: out<=0;
   23115: out<=0;
   23116: out<=0;
   23117: out<=1;
   23118: out<=1;
   23119: out<=0;
   23120: out<=0;
   23121: out<=0;
   23122: out<=1;
   23123: out<=1;
   23124: out<=1;
   23125: out<=0;
   23126: out<=1;
   23127: out<=0;
   23128: out<=0;
   23129: out<=1;
   23130: out<=1;
   23131: out<=0;
   23132: out<=1;
   23133: out<=1;
   23134: out<=1;
   23135: out<=1;
   23136: out<=0;
   23137: out<=0;
   23138: out<=0;
   23139: out<=0;
   23140: out<=1;
   23141: out<=0;
   23142: out<=0;
   23143: out<=1;
   23144: out<=1;
   23145: out<=0;
   23146: out<=1;
   23147: out<=0;
   23148: out<=0;
   23149: out<=0;
   23150: out<=1;
   23151: out<=1;
   23152: out<=1;
   23153: out<=0;
   23154: out<=0;
   23155: out<=1;
   23156: out<=1;
   23157: out<=1;
   23158: out<=1;
   23159: out<=1;
   23160: out<=1;
   23161: out<=1;
   23162: out<=0;
   23163: out<=0;
   23164: out<=1;
   23165: out<=0;
   23166: out<=1;
   23167: out<=0;
   23168: out<=0;
   23169: out<=1;
   23170: out<=0;
   23171: out<=1;
   23172: out<=0;
   23173: out<=0;
   23174: out<=1;
   23175: out<=1;
   23176: out<=1;
   23177: out<=1;
   23178: out<=1;
   23179: out<=1;
   23180: out<=1;
   23181: out<=0;
   23182: out<=0;
   23183: out<=1;
   23184: out<=1;
   23185: out<=1;
   23186: out<=0;
   23187: out<=0;
   23188: out<=0;
   23189: out<=1;
   23190: out<=0;
   23191: out<=1;
   23192: out<=1;
   23193: out<=0;
   23194: out<=0;
   23195: out<=1;
   23196: out<=0;
   23197: out<=0;
   23198: out<=0;
   23199: out<=0;
   23200: out<=0;
   23201: out<=0;
   23202: out<=0;
   23203: out<=0;
   23204: out<=1;
   23205: out<=0;
   23206: out<=0;
   23207: out<=1;
   23208: out<=1;
   23209: out<=0;
   23210: out<=1;
   23211: out<=0;
   23212: out<=0;
   23213: out<=0;
   23214: out<=1;
   23215: out<=1;
   23216: out<=1;
   23217: out<=0;
   23218: out<=0;
   23219: out<=1;
   23220: out<=1;
   23221: out<=1;
   23222: out<=1;
   23223: out<=1;
   23224: out<=1;
   23225: out<=1;
   23226: out<=0;
   23227: out<=0;
   23228: out<=1;
   23229: out<=0;
   23230: out<=1;
   23231: out<=0;
   23232: out<=0;
   23233: out<=1;
   23234: out<=0;
   23235: out<=1;
   23236: out<=0;
   23237: out<=0;
   23238: out<=1;
   23239: out<=1;
   23240: out<=1;
   23241: out<=1;
   23242: out<=1;
   23243: out<=1;
   23244: out<=1;
   23245: out<=0;
   23246: out<=0;
   23247: out<=1;
   23248: out<=0;
   23249: out<=0;
   23250: out<=1;
   23251: out<=1;
   23252: out<=1;
   23253: out<=0;
   23254: out<=1;
   23255: out<=0;
   23256: out<=0;
   23257: out<=1;
   23258: out<=1;
   23259: out<=0;
   23260: out<=1;
   23261: out<=1;
   23262: out<=1;
   23263: out<=1;
   23264: out<=1;
   23265: out<=1;
   23266: out<=1;
   23267: out<=1;
   23268: out<=0;
   23269: out<=1;
   23270: out<=1;
   23271: out<=0;
   23272: out<=0;
   23273: out<=1;
   23274: out<=0;
   23275: out<=1;
   23276: out<=1;
   23277: out<=1;
   23278: out<=0;
   23279: out<=0;
   23280: out<=1;
   23281: out<=0;
   23282: out<=0;
   23283: out<=1;
   23284: out<=1;
   23285: out<=1;
   23286: out<=1;
   23287: out<=1;
   23288: out<=1;
   23289: out<=1;
   23290: out<=0;
   23291: out<=0;
   23292: out<=1;
   23293: out<=0;
   23294: out<=1;
   23295: out<=0;
   23296: out<=0;
   23297: out<=0;
   23298: out<=1;
   23299: out<=1;
   23300: out<=1;
   23301: out<=0;
   23302: out<=1;
   23303: out<=0;
   23304: out<=0;
   23305: out<=1;
   23306: out<=1;
   23307: out<=0;
   23308: out<=1;
   23309: out<=1;
   23310: out<=1;
   23311: out<=1;
   23312: out<=1;
   23313: out<=0;
   23314: out<=1;
   23315: out<=0;
   23316: out<=1;
   23317: out<=1;
   23318: out<=0;
   23319: out<=0;
   23320: out<=0;
   23321: out<=0;
   23322: out<=0;
   23323: out<=0;
   23324: out<=0;
   23325: out<=1;
   23326: out<=1;
   23327: out<=0;
   23328: out<=1;
   23329: out<=0;
   23330: out<=0;
   23331: out<=1;
   23332: out<=1;
   23333: out<=1;
   23334: out<=1;
   23335: out<=1;
   23336: out<=1;
   23337: out<=1;
   23338: out<=0;
   23339: out<=0;
   23340: out<=1;
   23341: out<=0;
   23342: out<=1;
   23343: out<=0;
   23344: out<=0;
   23345: out<=0;
   23346: out<=0;
   23347: out<=0;
   23348: out<=1;
   23349: out<=0;
   23350: out<=0;
   23351: out<=1;
   23352: out<=1;
   23353: out<=0;
   23354: out<=1;
   23355: out<=0;
   23356: out<=0;
   23357: out<=0;
   23358: out<=1;
   23359: out<=1;
   23360: out<=1;
   23361: out<=1;
   23362: out<=0;
   23363: out<=0;
   23364: out<=0;
   23365: out<=1;
   23366: out<=0;
   23367: out<=1;
   23368: out<=1;
   23369: out<=0;
   23370: out<=0;
   23371: out<=1;
   23372: out<=0;
   23373: out<=0;
   23374: out<=0;
   23375: out<=0;
   23376: out<=1;
   23377: out<=0;
   23378: out<=1;
   23379: out<=0;
   23380: out<=1;
   23381: out<=1;
   23382: out<=0;
   23383: out<=0;
   23384: out<=0;
   23385: out<=0;
   23386: out<=0;
   23387: out<=0;
   23388: out<=0;
   23389: out<=1;
   23390: out<=1;
   23391: out<=0;
   23392: out<=1;
   23393: out<=0;
   23394: out<=0;
   23395: out<=1;
   23396: out<=1;
   23397: out<=1;
   23398: out<=1;
   23399: out<=1;
   23400: out<=1;
   23401: out<=1;
   23402: out<=0;
   23403: out<=0;
   23404: out<=1;
   23405: out<=0;
   23406: out<=1;
   23407: out<=0;
   23408: out<=1;
   23409: out<=1;
   23410: out<=1;
   23411: out<=1;
   23412: out<=0;
   23413: out<=1;
   23414: out<=1;
   23415: out<=0;
   23416: out<=0;
   23417: out<=1;
   23418: out<=0;
   23419: out<=1;
   23420: out<=1;
   23421: out<=1;
   23422: out<=0;
   23423: out<=0;
   23424: out<=0;
   23425: out<=0;
   23426: out<=1;
   23427: out<=1;
   23428: out<=1;
   23429: out<=0;
   23430: out<=1;
   23431: out<=0;
   23432: out<=0;
   23433: out<=1;
   23434: out<=1;
   23435: out<=0;
   23436: out<=1;
   23437: out<=1;
   23438: out<=1;
   23439: out<=1;
   23440: out<=0;
   23441: out<=1;
   23442: out<=0;
   23443: out<=1;
   23444: out<=0;
   23445: out<=0;
   23446: out<=1;
   23447: out<=1;
   23448: out<=1;
   23449: out<=1;
   23450: out<=1;
   23451: out<=1;
   23452: out<=1;
   23453: out<=0;
   23454: out<=0;
   23455: out<=1;
   23456: out<=1;
   23457: out<=0;
   23458: out<=0;
   23459: out<=1;
   23460: out<=1;
   23461: out<=1;
   23462: out<=1;
   23463: out<=1;
   23464: out<=1;
   23465: out<=1;
   23466: out<=0;
   23467: out<=0;
   23468: out<=1;
   23469: out<=0;
   23470: out<=1;
   23471: out<=0;
   23472: out<=1;
   23473: out<=1;
   23474: out<=1;
   23475: out<=1;
   23476: out<=0;
   23477: out<=1;
   23478: out<=1;
   23479: out<=0;
   23480: out<=0;
   23481: out<=1;
   23482: out<=0;
   23483: out<=1;
   23484: out<=1;
   23485: out<=1;
   23486: out<=0;
   23487: out<=0;
   23488: out<=1;
   23489: out<=1;
   23490: out<=0;
   23491: out<=0;
   23492: out<=0;
   23493: out<=1;
   23494: out<=0;
   23495: out<=1;
   23496: out<=1;
   23497: out<=0;
   23498: out<=0;
   23499: out<=1;
   23500: out<=0;
   23501: out<=0;
   23502: out<=0;
   23503: out<=0;
   23504: out<=0;
   23505: out<=1;
   23506: out<=0;
   23507: out<=1;
   23508: out<=0;
   23509: out<=0;
   23510: out<=1;
   23511: out<=1;
   23512: out<=1;
   23513: out<=1;
   23514: out<=1;
   23515: out<=1;
   23516: out<=1;
   23517: out<=0;
   23518: out<=0;
   23519: out<=1;
   23520: out<=1;
   23521: out<=0;
   23522: out<=0;
   23523: out<=1;
   23524: out<=1;
   23525: out<=1;
   23526: out<=1;
   23527: out<=1;
   23528: out<=1;
   23529: out<=1;
   23530: out<=0;
   23531: out<=0;
   23532: out<=1;
   23533: out<=0;
   23534: out<=1;
   23535: out<=0;
   23536: out<=0;
   23537: out<=0;
   23538: out<=0;
   23539: out<=0;
   23540: out<=1;
   23541: out<=0;
   23542: out<=0;
   23543: out<=1;
   23544: out<=1;
   23545: out<=0;
   23546: out<=1;
   23547: out<=0;
   23548: out<=0;
   23549: out<=0;
   23550: out<=1;
   23551: out<=1;
   23552: out<=0;
   23553: out<=1;
   23554: out<=1;
   23555: out<=0;
   23556: out<=1;
   23557: out<=1;
   23558: out<=1;
   23559: out<=1;
   23560: out<=1;
   23561: out<=1;
   23562: out<=0;
   23563: out<=0;
   23564: out<=0;
   23565: out<=1;
   23566: out<=0;
   23567: out<=1;
   23568: out<=1;
   23569: out<=1;
   23570: out<=1;
   23571: out<=1;
   23572: out<=1;
   23573: out<=0;
   23574: out<=0;
   23575: out<=1;
   23576: out<=1;
   23577: out<=0;
   23578: out<=1;
   23579: out<=0;
   23580: out<=1;
   23581: out<=1;
   23582: out<=0;
   23583: out<=0;
   23584: out<=0;
   23585: out<=0;
   23586: out<=1;
   23587: out<=1;
   23588: out<=0;
   23589: out<=1;
   23590: out<=0;
   23591: out<=1;
   23592: out<=1;
   23593: out<=0;
   23594: out<=0;
   23595: out<=1;
   23596: out<=1;
   23597: out<=1;
   23598: out<=1;
   23599: out<=1;
   23600: out<=1;
   23601: out<=0;
   23602: out<=1;
   23603: out<=0;
   23604: out<=0;
   23605: out<=0;
   23606: out<=1;
   23607: out<=1;
   23608: out<=1;
   23609: out<=1;
   23610: out<=1;
   23611: out<=1;
   23612: out<=0;
   23613: out<=1;
   23614: out<=1;
   23615: out<=0;
   23616: out<=0;
   23617: out<=1;
   23618: out<=1;
   23619: out<=0;
   23620: out<=1;
   23621: out<=1;
   23622: out<=1;
   23623: out<=1;
   23624: out<=1;
   23625: out<=1;
   23626: out<=0;
   23627: out<=0;
   23628: out<=0;
   23629: out<=1;
   23630: out<=0;
   23631: out<=1;
   23632: out<=0;
   23633: out<=0;
   23634: out<=0;
   23635: out<=0;
   23636: out<=0;
   23637: out<=1;
   23638: out<=1;
   23639: out<=0;
   23640: out<=0;
   23641: out<=1;
   23642: out<=0;
   23643: out<=1;
   23644: out<=0;
   23645: out<=0;
   23646: out<=1;
   23647: out<=1;
   23648: out<=1;
   23649: out<=1;
   23650: out<=0;
   23651: out<=0;
   23652: out<=1;
   23653: out<=0;
   23654: out<=1;
   23655: out<=0;
   23656: out<=0;
   23657: out<=1;
   23658: out<=1;
   23659: out<=0;
   23660: out<=0;
   23661: out<=0;
   23662: out<=0;
   23663: out<=0;
   23664: out<=1;
   23665: out<=0;
   23666: out<=1;
   23667: out<=0;
   23668: out<=0;
   23669: out<=0;
   23670: out<=1;
   23671: out<=1;
   23672: out<=1;
   23673: out<=1;
   23674: out<=1;
   23675: out<=1;
   23676: out<=0;
   23677: out<=1;
   23678: out<=1;
   23679: out<=0;
   23680: out<=0;
   23681: out<=1;
   23682: out<=1;
   23683: out<=0;
   23684: out<=1;
   23685: out<=1;
   23686: out<=1;
   23687: out<=1;
   23688: out<=1;
   23689: out<=1;
   23690: out<=0;
   23691: out<=0;
   23692: out<=0;
   23693: out<=1;
   23694: out<=0;
   23695: out<=1;
   23696: out<=0;
   23697: out<=0;
   23698: out<=0;
   23699: out<=0;
   23700: out<=0;
   23701: out<=1;
   23702: out<=1;
   23703: out<=0;
   23704: out<=0;
   23705: out<=1;
   23706: out<=0;
   23707: out<=1;
   23708: out<=0;
   23709: out<=0;
   23710: out<=1;
   23711: out<=1;
   23712: out<=0;
   23713: out<=0;
   23714: out<=1;
   23715: out<=1;
   23716: out<=0;
   23717: out<=1;
   23718: out<=0;
   23719: out<=1;
   23720: out<=1;
   23721: out<=0;
   23722: out<=0;
   23723: out<=1;
   23724: out<=1;
   23725: out<=1;
   23726: out<=1;
   23727: out<=1;
   23728: out<=0;
   23729: out<=1;
   23730: out<=0;
   23731: out<=1;
   23732: out<=1;
   23733: out<=1;
   23734: out<=0;
   23735: out<=0;
   23736: out<=0;
   23737: out<=0;
   23738: out<=0;
   23739: out<=0;
   23740: out<=1;
   23741: out<=0;
   23742: out<=0;
   23743: out<=1;
   23744: out<=0;
   23745: out<=1;
   23746: out<=1;
   23747: out<=0;
   23748: out<=1;
   23749: out<=1;
   23750: out<=1;
   23751: out<=1;
   23752: out<=1;
   23753: out<=1;
   23754: out<=0;
   23755: out<=0;
   23756: out<=0;
   23757: out<=1;
   23758: out<=0;
   23759: out<=1;
   23760: out<=1;
   23761: out<=1;
   23762: out<=1;
   23763: out<=1;
   23764: out<=1;
   23765: out<=0;
   23766: out<=0;
   23767: out<=1;
   23768: out<=1;
   23769: out<=0;
   23770: out<=1;
   23771: out<=0;
   23772: out<=1;
   23773: out<=1;
   23774: out<=0;
   23775: out<=0;
   23776: out<=1;
   23777: out<=1;
   23778: out<=0;
   23779: out<=0;
   23780: out<=1;
   23781: out<=0;
   23782: out<=1;
   23783: out<=0;
   23784: out<=0;
   23785: out<=1;
   23786: out<=1;
   23787: out<=0;
   23788: out<=0;
   23789: out<=0;
   23790: out<=0;
   23791: out<=0;
   23792: out<=0;
   23793: out<=1;
   23794: out<=0;
   23795: out<=1;
   23796: out<=1;
   23797: out<=1;
   23798: out<=0;
   23799: out<=0;
   23800: out<=0;
   23801: out<=0;
   23802: out<=0;
   23803: out<=0;
   23804: out<=1;
   23805: out<=0;
   23806: out<=0;
   23807: out<=1;
   23808: out<=0;
   23809: out<=0;
   23810: out<=0;
   23811: out<=0;
   23812: out<=0;
   23813: out<=1;
   23814: out<=1;
   23815: out<=0;
   23816: out<=0;
   23817: out<=1;
   23818: out<=0;
   23819: out<=1;
   23820: out<=0;
   23821: out<=0;
   23822: out<=1;
   23823: out<=1;
   23824: out<=0;
   23825: out<=1;
   23826: out<=1;
   23827: out<=0;
   23828: out<=1;
   23829: out<=1;
   23830: out<=1;
   23831: out<=1;
   23832: out<=1;
   23833: out<=1;
   23834: out<=0;
   23835: out<=0;
   23836: out<=0;
   23837: out<=1;
   23838: out<=0;
   23839: out<=1;
   23840: out<=1;
   23841: out<=0;
   23842: out<=1;
   23843: out<=0;
   23844: out<=0;
   23845: out<=0;
   23846: out<=1;
   23847: out<=1;
   23848: out<=1;
   23849: out<=1;
   23850: out<=1;
   23851: out<=1;
   23852: out<=0;
   23853: out<=1;
   23854: out<=1;
   23855: out<=0;
   23856: out<=1;
   23857: out<=1;
   23858: out<=0;
   23859: out<=0;
   23860: out<=1;
   23861: out<=0;
   23862: out<=1;
   23863: out<=0;
   23864: out<=0;
   23865: out<=1;
   23866: out<=1;
   23867: out<=0;
   23868: out<=0;
   23869: out<=0;
   23870: out<=0;
   23871: out<=0;
   23872: out<=1;
   23873: out<=1;
   23874: out<=1;
   23875: out<=1;
   23876: out<=1;
   23877: out<=0;
   23878: out<=0;
   23879: out<=1;
   23880: out<=1;
   23881: out<=0;
   23882: out<=1;
   23883: out<=0;
   23884: out<=1;
   23885: out<=1;
   23886: out<=0;
   23887: out<=0;
   23888: out<=0;
   23889: out<=1;
   23890: out<=1;
   23891: out<=0;
   23892: out<=1;
   23893: out<=1;
   23894: out<=1;
   23895: out<=1;
   23896: out<=1;
   23897: out<=1;
   23898: out<=0;
   23899: out<=0;
   23900: out<=0;
   23901: out<=1;
   23902: out<=0;
   23903: out<=1;
   23904: out<=1;
   23905: out<=0;
   23906: out<=1;
   23907: out<=0;
   23908: out<=0;
   23909: out<=0;
   23910: out<=1;
   23911: out<=1;
   23912: out<=1;
   23913: out<=1;
   23914: out<=1;
   23915: out<=1;
   23916: out<=0;
   23917: out<=1;
   23918: out<=1;
   23919: out<=0;
   23920: out<=0;
   23921: out<=0;
   23922: out<=1;
   23923: out<=1;
   23924: out<=0;
   23925: out<=1;
   23926: out<=0;
   23927: out<=1;
   23928: out<=1;
   23929: out<=0;
   23930: out<=0;
   23931: out<=1;
   23932: out<=1;
   23933: out<=1;
   23934: out<=1;
   23935: out<=1;
   23936: out<=1;
   23937: out<=1;
   23938: out<=1;
   23939: out<=1;
   23940: out<=1;
   23941: out<=0;
   23942: out<=0;
   23943: out<=1;
   23944: out<=1;
   23945: out<=0;
   23946: out<=1;
   23947: out<=0;
   23948: out<=1;
   23949: out<=1;
   23950: out<=0;
   23951: out<=0;
   23952: out<=0;
   23953: out<=1;
   23954: out<=1;
   23955: out<=0;
   23956: out<=1;
   23957: out<=1;
   23958: out<=1;
   23959: out<=1;
   23960: out<=1;
   23961: out<=1;
   23962: out<=0;
   23963: out<=0;
   23964: out<=0;
   23965: out<=1;
   23966: out<=0;
   23967: out<=1;
   23968: out<=0;
   23969: out<=1;
   23970: out<=0;
   23971: out<=1;
   23972: out<=1;
   23973: out<=1;
   23974: out<=0;
   23975: out<=0;
   23976: out<=0;
   23977: out<=0;
   23978: out<=0;
   23979: out<=0;
   23980: out<=1;
   23981: out<=0;
   23982: out<=0;
   23983: out<=1;
   23984: out<=1;
   23985: out<=1;
   23986: out<=0;
   23987: out<=0;
   23988: out<=1;
   23989: out<=0;
   23990: out<=1;
   23991: out<=0;
   23992: out<=0;
   23993: out<=1;
   23994: out<=1;
   23995: out<=0;
   23996: out<=0;
   23997: out<=0;
   23998: out<=0;
   23999: out<=0;
   24000: out<=0;
   24001: out<=0;
   24002: out<=0;
   24003: out<=0;
   24004: out<=0;
   24005: out<=1;
   24006: out<=1;
   24007: out<=0;
   24008: out<=0;
   24009: out<=1;
   24010: out<=0;
   24011: out<=1;
   24012: out<=0;
   24013: out<=0;
   24014: out<=1;
   24015: out<=1;
   24016: out<=0;
   24017: out<=1;
   24018: out<=1;
   24019: out<=0;
   24020: out<=1;
   24021: out<=1;
   24022: out<=1;
   24023: out<=1;
   24024: out<=1;
   24025: out<=1;
   24026: out<=0;
   24027: out<=0;
   24028: out<=0;
   24029: out<=1;
   24030: out<=0;
   24031: out<=1;
   24032: out<=0;
   24033: out<=1;
   24034: out<=0;
   24035: out<=1;
   24036: out<=1;
   24037: out<=1;
   24038: out<=0;
   24039: out<=0;
   24040: out<=0;
   24041: out<=0;
   24042: out<=0;
   24043: out<=0;
   24044: out<=1;
   24045: out<=0;
   24046: out<=0;
   24047: out<=1;
   24048: out<=0;
   24049: out<=0;
   24050: out<=1;
   24051: out<=1;
   24052: out<=0;
   24053: out<=1;
   24054: out<=0;
   24055: out<=1;
   24056: out<=1;
   24057: out<=0;
   24058: out<=0;
   24059: out<=1;
   24060: out<=1;
   24061: out<=1;
   24062: out<=1;
   24063: out<=1;
   24064: out<=0;
   24065: out<=0;
   24066: out<=1;
   24067: out<=1;
   24068: out<=0;
   24069: out<=1;
   24070: out<=0;
   24071: out<=1;
   24072: out<=1;
   24073: out<=0;
   24074: out<=0;
   24075: out<=1;
   24076: out<=1;
   24077: out<=1;
   24078: out<=1;
   24079: out<=1;
   24080: out<=0;
   24081: out<=1;
   24082: out<=0;
   24083: out<=1;
   24084: out<=1;
   24085: out<=1;
   24086: out<=0;
   24087: out<=0;
   24088: out<=0;
   24089: out<=0;
   24090: out<=0;
   24091: out<=0;
   24092: out<=1;
   24093: out<=0;
   24094: out<=0;
   24095: out<=1;
   24096: out<=0;
   24097: out<=1;
   24098: out<=1;
   24099: out<=0;
   24100: out<=1;
   24101: out<=1;
   24102: out<=1;
   24103: out<=1;
   24104: out<=1;
   24105: out<=1;
   24106: out<=0;
   24107: out<=0;
   24108: out<=0;
   24109: out<=1;
   24110: out<=0;
   24111: out<=1;
   24112: out<=0;
   24113: out<=0;
   24114: out<=0;
   24115: out<=0;
   24116: out<=0;
   24117: out<=1;
   24118: out<=1;
   24119: out<=0;
   24120: out<=0;
   24121: out<=1;
   24122: out<=0;
   24123: out<=1;
   24124: out<=0;
   24125: out<=0;
   24126: out<=1;
   24127: out<=1;
   24128: out<=1;
   24129: out<=1;
   24130: out<=0;
   24131: out<=0;
   24132: out<=1;
   24133: out<=0;
   24134: out<=1;
   24135: out<=0;
   24136: out<=0;
   24137: out<=1;
   24138: out<=1;
   24139: out<=0;
   24140: out<=0;
   24141: out<=0;
   24142: out<=0;
   24143: out<=0;
   24144: out<=0;
   24145: out<=1;
   24146: out<=0;
   24147: out<=1;
   24148: out<=1;
   24149: out<=1;
   24150: out<=0;
   24151: out<=0;
   24152: out<=0;
   24153: out<=0;
   24154: out<=0;
   24155: out<=0;
   24156: out<=1;
   24157: out<=0;
   24158: out<=0;
   24159: out<=1;
   24160: out<=0;
   24161: out<=1;
   24162: out<=1;
   24163: out<=0;
   24164: out<=1;
   24165: out<=1;
   24166: out<=1;
   24167: out<=1;
   24168: out<=1;
   24169: out<=1;
   24170: out<=0;
   24171: out<=0;
   24172: out<=0;
   24173: out<=1;
   24174: out<=0;
   24175: out<=1;
   24176: out<=1;
   24177: out<=1;
   24178: out<=1;
   24179: out<=1;
   24180: out<=1;
   24181: out<=0;
   24182: out<=0;
   24183: out<=1;
   24184: out<=1;
   24185: out<=0;
   24186: out<=1;
   24187: out<=0;
   24188: out<=1;
   24189: out<=1;
   24190: out<=0;
   24191: out<=0;
   24192: out<=0;
   24193: out<=0;
   24194: out<=1;
   24195: out<=1;
   24196: out<=0;
   24197: out<=1;
   24198: out<=0;
   24199: out<=1;
   24200: out<=1;
   24201: out<=0;
   24202: out<=0;
   24203: out<=1;
   24204: out<=1;
   24205: out<=1;
   24206: out<=1;
   24207: out<=1;
   24208: out<=1;
   24209: out<=0;
   24210: out<=1;
   24211: out<=0;
   24212: out<=0;
   24213: out<=0;
   24214: out<=1;
   24215: out<=1;
   24216: out<=1;
   24217: out<=1;
   24218: out<=1;
   24219: out<=1;
   24220: out<=0;
   24221: out<=1;
   24222: out<=1;
   24223: out<=0;
   24224: out<=0;
   24225: out<=1;
   24226: out<=1;
   24227: out<=0;
   24228: out<=1;
   24229: out<=1;
   24230: out<=1;
   24231: out<=1;
   24232: out<=1;
   24233: out<=1;
   24234: out<=0;
   24235: out<=0;
   24236: out<=0;
   24237: out<=1;
   24238: out<=0;
   24239: out<=1;
   24240: out<=1;
   24241: out<=1;
   24242: out<=1;
   24243: out<=1;
   24244: out<=1;
   24245: out<=0;
   24246: out<=0;
   24247: out<=1;
   24248: out<=1;
   24249: out<=0;
   24250: out<=1;
   24251: out<=0;
   24252: out<=1;
   24253: out<=1;
   24254: out<=0;
   24255: out<=0;
   24256: out<=1;
   24257: out<=1;
   24258: out<=0;
   24259: out<=0;
   24260: out<=1;
   24261: out<=0;
   24262: out<=1;
   24263: out<=0;
   24264: out<=0;
   24265: out<=1;
   24266: out<=1;
   24267: out<=0;
   24268: out<=0;
   24269: out<=0;
   24270: out<=0;
   24271: out<=0;
   24272: out<=1;
   24273: out<=0;
   24274: out<=1;
   24275: out<=0;
   24276: out<=0;
   24277: out<=0;
   24278: out<=1;
   24279: out<=1;
   24280: out<=1;
   24281: out<=1;
   24282: out<=1;
   24283: out<=1;
   24284: out<=0;
   24285: out<=1;
   24286: out<=1;
   24287: out<=0;
   24288: out<=0;
   24289: out<=1;
   24290: out<=1;
   24291: out<=0;
   24292: out<=1;
   24293: out<=1;
   24294: out<=1;
   24295: out<=1;
   24296: out<=1;
   24297: out<=1;
   24298: out<=0;
   24299: out<=0;
   24300: out<=0;
   24301: out<=1;
   24302: out<=0;
   24303: out<=1;
   24304: out<=0;
   24305: out<=0;
   24306: out<=0;
   24307: out<=0;
   24308: out<=0;
   24309: out<=1;
   24310: out<=1;
   24311: out<=0;
   24312: out<=0;
   24313: out<=1;
   24314: out<=0;
   24315: out<=1;
   24316: out<=0;
   24317: out<=0;
   24318: out<=1;
   24319: out<=1;
   24320: out<=0;
   24321: out<=1;
   24322: out<=0;
   24323: out<=1;
   24324: out<=1;
   24325: out<=1;
   24326: out<=0;
   24327: out<=0;
   24328: out<=0;
   24329: out<=0;
   24330: out<=0;
   24331: out<=0;
   24332: out<=1;
   24333: out<=0;
   24334: out<=0;
   24335: out<=1;
   24336: out<=1;
   24337: out<=1;
   24338: out<=0;
   24339: out<=0;
   24340: out<=1;
   24341: out<=0;
   24342: out<=1;
   24343: out<=0;
   24344: out<=0;
   24345: out<=1;
   24346: out<=1;
   24347: out<=0;
   24348: out<=0;
   24349: out<=0;
   24350: out<=0;
   24351: out<=0;
   24352: out<=1;
   24353: out<=1;
   24354: out<=1;
   24355: out<=1;
   24356: out<=1;
   24357: out<=0;
   24358: out<=0;
   24359: out<=1;
   24360: out<=1;
   24361: out<=0;
   24362: out<=1;
   24363: out<=0;
   24364: out<=1;
   24365: out<=1;
   24366: out<=0;
   24367: out<=0;
   24368: out<=0;
   24369: out<=1;
   24370: out<=1;
   24371: out<=0;
   24372: out<=1;
   24373: out<=1;
   24374: out<=1;
   24375: out<=1;
   24376: out<=1;
   24377: out<=1;
   24378: out<=0;
   24379: out<=0;
   24380: out<=0;
   24381: out<=1;
   24382: out<=0;
   24383: out<=1;
   24384: out<=0;
   24385: out<=1;
   24386: out<=0;
   24387: out<=1;
   24388: out<=1;
   24389: out<=1;
   24390: out<=0;
   24391: out<=0;
   24392: out<=0;
   24393: out<=0;
   24394: out<=0;
   24395: out<=0;
   24396: out<=1;
   24397: out<=0;
   24398: out<=0;
   24399: out<=1;
   24400: out<=0;
   24401: out<=0;
   24402: out<=1;
   24403: out<=1;
   24404: out<=0;
   24405: out<=1;
   24406: out<=0;
   24407: out<=1;
   24408: out<=1;
   24409: out<=0;
   24410: out<=0;
   24411: out<=1;
   24412: out<=1;
   24413: out<=1;
   24414: out<=1;
   24415: out<=1;
   24416: out<=0;
   24417: out<=0;
   24418: out<=0;
   24419: out<=0;
   24420: out<=0;
   24421: out<=1;
   24422: out<=1;
   24423: out<=0;
   24424: out<=0;
   24425: out<=1;
   24426: out<=0;
   24427: out<=1;
   24428: out<=0;
   24429: out<=0;
   24430: out<=1;
   24431: out<=1;
   24432: out<=0;
   24433: out<=1;
   24434: out<=1;
   24435: out<=0;
   24436: out<=1;
   24437: out<=1;
   24438: out<=1;
   24439: out<=1;
   24440: out<=1;
   24441: out<=1;
   24442: out<=0;
   24443: out<=0;
   24444: out<=0;
   24445: out<=1;
   24446: out<=0;
   24447: out<=1;
   24448: out<=1;
   24449: out<=0;
   24450: out<=1;
   24451: out<=0;
   24452: out<=0;
   24453: out<=0;
   24454: out<=1;
   24455: out<=1;
   24456: out<=1;
   24457: out<=1;
   24458: out<=1;
   24459: out<=1;
   24460: out<=0;
   24461: out<=1;
   24462: out<=1;
   24463: out<=0;
   24464: out<=1;
   24465: out<=1;
   24466: out<=0;
   24467: out<=0;
   24468: out<=1;
   24469: out<=0;
   24470: out<=1;
   24471: out<=0;
   24472: out<=0;
   24473: out<=1;
   24474: out<=1;
   24475: out<=0;
   24476: out<=0;
   24477: out<=0;
   24478: out<=0;
   24479: out<=0;
   24480: out<=0;
   24481: out<=0;
   24482: out<=0;
   24483: out<=0;
   24484: out<=0;
   24485: out<=1;
   24486: out<=1;
   24487: out<=0;
   24488: out<=0;
   24489: out<=1;
   24490: out<=0;
   24491: out<=1;
   24492: out<=0;
   24493: out<=0;
   24494: out<=1;
   24495: out<=1;
   24496: out<=0;
   24497: out<=1;
   24498: out<=1;
   24499: out<=0;
   24500: out<=1;
   24501: out<=1;
   24502: out<=1;
   24503: out<=1;
   24504: out<=1;
   24505: out<=1;
   24506: out<=0;
   24507: out<=0;
   24508: out<=0;
   24509: out<=1;
   24510: out<=0;
   24511: out<=1;
   24512: out<=1;
   24513: out<=0;
   24514: out<=1;
   24515: out<=0;
   24516: out<=0;
   24517: out<=0;
   24518: out<=1;
   24519: out<=1;
   24520: out<=1;
   24521: out<=1;
   24522: out<=1;
   24523: out<=1;
   24524: out<=0;
   24525: out<=1;
   24526: out<=1;
   24527: out<=0;
   24528: out<=0;
   24529: out<=0;
   24530: out<=1;
   24531: out<=1;
   24532: out<=0;
   24533: out<=1;
   24534: out<=0;
   24535: out<=1;
   24536: out<=1;
   24537: out<=0;
   24538: out<=0;
   24539: out<=1;
   24540: out<=1;
   24541: out<=1;
   24542: out<=1;
   24543: out<=1;
   24544: out<=1;
   24545: out<=1;
   24546: out<=1;
   24547: out<=1;
   24548: out<=1;
   24549: out<=0;
   24550: out<=0;
   24551: out<=1;
   24552: out<=1;
   24553: out<=0;
   24554: out<=1;
   24555: out<=0;
   24556: out<=1;
   24557: out<=1;
   24558: out<=0;
   24559: out<=0;
   24560: out<=0;
   24561: out<=1;
   24562: out<=1;
   24563: out<=0;
   24564: out<=1;
   24565: out<=1;
   24566: out<=1;
   24567: out<=1;
   24568: out<=1;
   24569: out<=1;
   24570: out<=0;
   24571: out<=0;
   24572: out<=0;
   24573: out<=1;
   24574: out<=0;
   24575: out<=1;
   24576: out<=0;
   24577: out<=1;
   24578: out<=0;
   24579: out<=1;
   24580: out<=1;
   24581: out<=1;
   24582: out<=0;
   24583: out<=0;
   24584: out<=0;
   24585: out<=0;
   24586: out<=0;
   24587: out<=0;
   24588: out<=1;
   24589: out<=0;
   24590: out<=0;
   24591: out<=1;
   24592: out<=1;
   24593: out<=1;
   24594: out<=0;
   24595: out<=0;
   24596: out<=1;
   24597: out<=0;
   24598: out<=1;
   24599: out<=0;
   24600: out<=0;
   24601: out<=1;
   24602: out<=1;
   24603: out<=0;
   24604: out<=0;
   24605: out<=0;
   24606: out<=0;
   24607: out<=0;
   24608: out<=0;
   24609: out<=0;
   24610: out<=0;
   24611: out<=0;
   24612: out<=0;
   24613: out<=1;
   24614: out<=1;
   24615: out<=0;
   24616: out<=0;
   24617: out<=1;
   24618: out<=0;
   24619: out<=1;
   24620: out<=0;
   24621: out<=0;
   24622: out<=1;
   24623: out<=1;
   24624: out<=1;
   24625: out<=0;
   24626: out<=0;
   24627: out<=1;
   24628: out<=0;
   24629: out<=0;
   24630: out<=0;
   24631: out<=0;
   24632: out<=0;
   24633: out<=0;
   24634: out<=1;
   24635: out<=1;
   24636: out<=1;
   24637: out<=0;
   24638: out<=1;
   24639: out<=0;
   24640: out<=0;
   24641: out<=1;
   24642: out<=0;
   24643: out<=1;
   24644: out<=1;
   24645: out<=1;
   24646: out<=0;
   24647: out<=0;
   24648: out<=0;
   24649: out<=0;
   24650: out<=0;
   24651: out<=0;
   24652: out<=1;
   24653: out<=0;
   24654: out<=0;
   24655: out<=1;
   24656: out<=0;
   24657: out<=0;
   24658: out<=1;
   24659: out<=1;
   24660: out<=0;
   24661: out<=1;
   24662: out<=0;
   24663: out<=1;
   24664: out<=1;
   24665: out<=0;
   24666: out<=0;
   24667: out<=1;
   24668: out<=1;
   24669: out<=1;
   24670: out<=1;
   24671: out<=1;
   24672: out<=1;
   24673: out<=1;
   24674: out<=1;
   24675: out<=1;
   24676: out<=1;
   24677: out<=0;
   24678: out<=0;
   24679: out<=1;
   24680: out<=1;
   24681: out<=0;
   24682: out<=1;
   24683: out<=0;
   24684: out<=1;
   24685: out<=1;
   24686: out<=0;
   24687: out<=0;
   24688: out<=1;
   24689: out<=0;
   24690: out<=0;
   24691: out<=1;
   24692: out<=0;
   24693: out<=0;
   24694: out<=0;
   24695: out<=0;
   24696: out<=0;
   24697: out<=0;
   24698: out<=1;
   24699: out<=1;
   24700: out<=1;
   24701: out<=0;
   24702: out<=1;
   24703: out<=0;
   24704: out<=1;
   24705: out<=0;
   24706: out<=1;
   24707: out<=0;
   24708: out<=0;
   24709: out<=0;
   24710: out<=1;
   24711: out<=1;
   24712: out<=1;
   24713: out<=1;
   24714: out<=1;
   24715: out<=1;
   24716: out<=0;
   24717: out<=1;
   24718: out<=1;
   24719: out<=0;
   24720: out<=1;
   24721: out<=1;
   24722: out<=0;
   24723: out<=0;
   24724: out<=1;
   24725: out<=0;
   24726: out<=1;
   24727: out<=0;
   24728: out<=0;
   24729: out<=1;
   24730: out<=1;
   24731: out<=0;
   24732: out<=0;
   24733: out<=0;
   24734: out<=0;
   24735: out<=0;
   24736: out<=1;
   24737: out<=1;
   24738: out<=1;
   24739: out<=1;
   24740: out<=1;
   24741: out<=0;
   24742: out<=0;
   24743: out<=1;
   24744: out<=1;
   24745: out<=0;
   24746: out<=1;
   24747: out<=0;
   24748: out<=1;
   24749: out<=1;
   24750: out<=0;
   24751: out<=0;
   24752: out<=1;
   24753: out<=0;
   24754: out<=0;
   24755: out<=1;
   24756: out<=0;
   24757: out<=0;
   24758: out<=0;
   24759: out<=0;
   24760: out<=0;
   24761: out<=0;
   24762: out<=1;
   24763: out<=1;
   24764: out<=1;
   24765: out<=0;
   24766: out<=1;
   24767: out<=0;
   24768: out<=1;
   24769: out<=0;
   24770: out<=1;
   24771: out<=0;
   24772: out<=0;
   24773: out<=0;
   24774: out<=1;
   24775: out<=1;
   24776: out<=1;
   24777: out<=1;
   24778: out<=1;
   24779: out<=1;
   24780: out<=0;
   24781: out<=1;
   24782: out<=1;
   24783: out<=0;
   24784: out<=0;
   24785: out<=0;
   24786: out<=1;
   24787: out<=1;
   24788: out<=0;
   24789: out<=1;
   24790: out<=0;
   24791: out<=1;
   24792: out<=1;
   24793: out<=0;
   24794: out<=0;
   24795: out<=1;
   24796: out<=1;
   24797: out<=1;
   24798: out<=1;
   24799: out<=1;
   24800: out<=0;
   24801: out<=0;
   24802: out<=0;
   24803: out<=0;
   24804: out<=0;
   24805: out<=1;
   24806: out<=1;
   24807: out<=0;
   24808: out<=0;
   24809: out<=1;
   24810: out<=0;
   24811: out<=1;
   24812: out<=0;
   24813: out<=0;
   24814: out<=1;
   24815: out<=1;
   24816: out<=1;
   24817: out<=0;
   24818: out<=0;
   24819: out<=1;
   24820: out<=0;
   24821: out<=0;
   24822: out<=0;
   24823: out<=0;
   24824: out<=0;
   24825: out<=0;
   24826: out<=1;
   24827: out<=1;
   24828: out<=1;
   24829: out<=0;
   24830: out<=1;
   24831: out<=0;
   24832: out<=0;
   24833: out<=0;
   24834: out<=1;
   24835: out<=1;
   24836: out<=0;
   24837: out<=1;
   24838: out<=0;
   24839: out<=1;
   24840: out<=1;
   24841: out<=0;
   24842: out<=0;
   24843: out<=1;
   24844: out<=1;
   24845: out<=1;
   24846: out<=1;
   24847: out<=1;
   24848: out<=0;
   24849: out<=1;
   24850: out<=0;
   24851: out<=1;
   24852: out<=1;
   24853: out<=1;
   24854: out<=0;
   24855: out<=0;
   24856: out<=0;
   24857: out<=0;
   24858: out<=0;
   24859: out<=0;
   24860: out<=1;
   24861: out<=0;
   24862: out<=0;
   24863: out<=1;
   24864: out<=1;
   24865: out<=0;
   24866: out<=0;
   24867: out<=1;
   24868: out<=0;
   24869: out<=0;
   24870: out<=0;
   24871: out<=0;
   24872: out<=0;
   24873: out<=0;
   24874: out<=1;
   24875: out<=1;
   24876: out<=1;
   24877: out<=0;
   24878: out<=1;
   24879: out<=0;
   24880: out<=1;
   24881: out<=1;
   24882: out<=1;
   24883: out<=1;
   24884: out<=1;
   24885: out<=0;
   24886: out<=0;
   24887: out<=1;
   24888: out<=1;
   24889: out<=0;
   24890: out<=1;
   24891: out<=0;
   24892: out<=1;
   24893: out<=1;
   24894: out<=0;
   24895: out<=0;
   24896: out<=1;
   24897: out<=1;
   24898: out<=0;
   24899: out<=0;
   24900: out<=1;
   24901: out<=0;
   24902: out<=1;
   24903: out<=0;
   24904: out<=0;
   24905: out<=1;
   24906: out<=1;
   24907: out<=0;
   24908: out<=0;
   24909: out<=0;
   24910: out<=0;
   24911: out<=0;
   24912: out<=0;
   24913: out<=1;
   24914: out<=0;
   24915: out<=1;
   24916: out<=1;
   24917: out<=1;
   24918: out<=0;
   24919: out<=0;
   24920: out<=0;
   24921: out<=0;
   24922: out<=0;
   24923: out<=0;
   24924: out<=1;
   24925: out<=0;
   24926: out<=0;
   24927: out<=1;
   24928: out<=1;
   24929: out<=0;
   24930: out<=0;
   24931: out<=1;
   24932: out<=0;
   24933: out<=0;
   24934: out<=0;
   24935: out<=0;
   24936: out<=0;
   24937: out<=0;
   24938: out<=1;
   24939: out<=1;
   24940: out<=1;
   24941: out<=0;
   24942: out<=1;
   24943: out<=0;
   24944: out<=0;
   24945: out<=0;
   24946: out<=0;
   24947: out<=0;
   24948: out<=0;
   24949: out<=1;
   24950: out<=1;
   24951: out<=0;
   24952: out<=0;
   24953: out<=1;
   24954: out<=0;
   24955: out<=1;
   24956: out<=0;
   24957: out<=0;
   24958: out<=1;
   24959: out<=1;
   24960: out<=0;
   24961: out<=0;
   24962: out<=1;
   24963: out<=1;
   24964: out<=0;
   24965: out<=1;
   24966: out<=0;
   24967: out<=1;
   24968: out<=1;
   24969: out<=0;
   24970: out<=0;
   24971: out<=1;
   24972: out<=1;
   24973: out<=1;
   24974: out<=1;
   24975: out<=1;
   24976: out<=1;
   24977: out<=0;
   24978: out<=1;
   24979: out<=0;
   24980: out<=0;
   24981: out<=0;
   24982: out<=1;
   24983: out<=1;
   24984: out<=1;
   24985: out<=1;
   24986: out<=1;
   24987: out<=1;
   24988: out<=0;
   24989: out<=1;
   24990: out<=1;
   24991: out<=0;
   24992: out<=1;
   24993: out<=0;
   24994: out<=0;
   24995: out<=1;
   24996: out<=0;
   24997: out<=0;
   24998: out<=0;
   24999: out<=0;
   25000: out<=0;
   25001: out<=0;
   25002: out<=1;
   25003: out<=1;
   25004: out<=1;
   25005: out<=0;
   25006: out<=1;
   25007: out<=0;
   25008: out<=0;
   25009: out<=0;
   25010: out<=0;
   25011: out<=0;
   25012: out<=0;
   25013: out<=1;
   25014: out<=1;
   25015: out<=0;
   25016: out<=0;
   25017: out<=1;
   25018: out<=0;
   25019: out<=1;
   25020: out<=0;
   25021: out<=0;
   25022: out<=1;
   25023: out<=1;
   25024: out<=1;
   25025: out<=1;
   25026: out<=0;
   25027: out<=0;
   25028: out<=1;
   25029: out<=0;
   25030: out<=1;
   25031: out<=0;
   25032: out<=0;
   25033: out<=1;
   25034: out<=1;
   25035: out<=0;
   25036: out<=0;
   25037: out<=0;
   25038: out<=0;
   25039: out<=0;
   25040: out<=1;
   25041: out<=0;
   25042: out<=1;
   25043: out<=0;
   25044: out<=0;
   25045: out<=0;
   25046: out<=1;
   25047: out<=1;
   25048: out<=1;
   25049: out<=1;
   25050: out<=1;
   25051: out<=1;
   25052: out<=0;
   25053: out<=1;
   25054: out<=1;
   25055: out<=0;
   25056: out<=1;
   25057: out<=0;
   25058: out<=0;
   25059: out<=1;
   25060: out<=0;
   25061: out<=0;
   25062: out<=0;
   25063: out<=0;
   25064: out<=0;
   25065: out<=0;
   25066: out<=1;
   25067: out<=1;
   25068: out<=1;
   25069: out<=0;
   25070: out<=1;
   25071: out<=0;
   25072: out<=1;
   25073: out<=1;
   25074: out<=1;
   25075: out<=1;
   25076: out<=1;
   25077: out<=0;
   25078: out<=0;
   25079: out<=1;
   25080: out<=1;
   25081: out<=0;
   25082: out<=1;
   25083: out<=0;
   25084: out<=1;
   25085: out<=1;
   25086: out<=0;
   25087: out<=0;
   25088: out<=1;
   25089: out<=1;
   25090: out<=1;
   25091: out<=1;
   25092: out<=1;
   25093: out<=0;
   25094: out<=0;
   25095: out<=1;
   25096: out<=1;
   25097: out<=0;
   25098: out<=1;
   25099: out<=0;
   25100: out<=1;
   25101: out<=1;
   25102: out<=0;
   25103: out<=0;
   25104: out<=1;
   25105: out<=0;
   25106: out<=0;
   25107: out<=1;
   25108: out<=0;
   25109: out<=0;
   25110: out<=0;
   25111: out<=0;
   25112: out<=0;
   25113: out<=0;
   25114: out<=1;
   25115: out<=1;
   25116: out<=1;
   25117: out<=0;
   25118: out<=1;
   25119: out<=0;
   25120: out<=1;
   25121: out<=0;
   25122: out<=1;
   25123: out<=0;
   25124: out<=0;
   25125: out<=0;
   25126: out<=1;
   25127: out<=1;
   25128: out<=1;
   25129: out<=1;
   25130: out<=1;
   25131: out<=1;
   25132: out<=0;
   25133: out<=1;
   25134: out<=1;
   25135: out<=0;
   25136: out<=1;
   25137: out<=1;
   25138: out<=0;
   25139: out<=0;
   25140: out<=1;
   25141: out<=0;
   25142: out<=1;
   25143: out<=0;
   25144: out<=0;
   25145: out<=1;
   25146: out<=1;
   25147: out<=0;
   25148: out<=0;
   25149: out<=0;
   25150: out<=0;
   25151: out<=0;
   25152: out<=0;
   25153: out<=0;
   25154: out<=0;
   25155: out<=0;
   25156: out<=0;
   25157: out<=1;
   25158: out<=1;
   25159: out<=0;
   25160: out<=0;
   25161: out<=1;
   25162: out<=0;
   25163: out<=1;
   25164: out<=0;
   25165: out<=0;
   25166: out<=1;
   25167: out<=1;
   25168: out<=1;
   25169: out<=0;
   25170: out<=0;
   25171: out<=1;
   25172: out<=0;
   25173: out<=0;
   25174: out<=0;
   25175: out<=0;
   25176: out<=0;
   25177: out<=0;
   25178: out<=1;
   25179: out<=1;
   25180: out<=1;
   25181: out<=0;
   25182: out<=1;
   25183: out<=0;
   25184: out<=1;
   25185: out<=0;
   25186: out<=1;
   25187: out<=0;
   25188: out<=0;
   25189: out<=0;
   25190: out<=1;
   25191: out<=1;
   25192: out<=1;
   25193: out<=1;
   25194: out<=1;
   25195: out<=1;
   25196: out<=0;
   25197: out<=1;
   25198: out<=1;
   25199: out<=0;
   25200: out<=0;
   25201: out<=0;
   25202: out<=1;
   25203: out<=1;
   25204: out<=0;
   25205: out<=1;
   25206: out<=0;
   25207: out<=1;
   25208: out<=1;
   25209: out<=0;
   25210: out<=0;
   25211: out<=1;
   25212: out<=1;
   25213: out<=1;
   25214: out<=1;
   25215: out<=1;
   25216: out<=0;
   25217: out<=0;
   25218: out<=0;
   25219: out<=0;
   25220: out<=0;
   25221: out<=1;
   25222: out<=1;
   25223: out<=0;
   25224: out<=0;
   25225: out<=1;
   25226: out<=0;
   25227: out<=1;
   25228: out<=0;
   25229: out<=0;
   25230: out<=1;
   25231: out<=1;
   25232: out<=1;
   25233: out<=0;
   25234: out<=0;
   25235: out<=1;
   25236: out<=0;
   25237: out<=0;
   25238: out<=0;
   25239: out<=0;
   25240: out<=0;
   25241: out<=0;
   25242: out<=1;
   25243: out<=1;
   25244: out<=1;
   25245: out<=0;
   25246: out<=1;
   25247: out<=0;
   25248: out<=0;
   25249: out<=1;
   25250: out<=0;
   25251: out<=1;
   25252: out<=1;
   25253: out<=1;
   25254: out<=0;
   25255: out<=0;
   25256: out<=0;
   25257: out<=0;
   25258: out<=0;
   25259: out<=0;
   25260: out<=1;
   25261: out<=0;
   25262: out<=0;
   25263: out<=1;
   25264: out<=1;
   25265: out<=1;
   25266: out<=0;
   25267: out<=0;
   25268: out<=1;
   25269: out<=0;
   25270: out<=1;
   25271: out<=0;
   25272: out<=0;
   25273: out<=1;
   25274: out<=1;
   25275: out<=0;
   25276: out<=0;
   25277: out<=0;
   25278: out<=0;
   25279: out<=0;
   25280: out<=1;
   25281: out<=1;
   25282: out<=1;
   25283: out<=1;
   25284: out<=1;
   25285: out<=0;
   25286: out<=0;
   25287: out<=1;
   25288: out<=1;
   25289: out<=0;
   25290: out<=1;
   25291: out<=0;
   25292: out<=1;
   25293: out<=1;
   25294: out<=0;
   25295: out<=0;
   25296: out<=1;
   25297: out<=0;
   25298: out<=0;
   25299: out<=1;
   25300: out<=0;
   25301: out<=0;
   25302: out<=0;
   25303: out<=0;
   25304: out<=0;
   25305: out<=0;
   25306: out<=1;
   25307: out<=1;
   25308: out<=1;
   25309: out<=0;
   25310: out<=1;
   25311: out<=0;
   25312: out<=0;
   25313: out<=1;
   25314: out<=0;
   25315: out<=1;
   25316: out<=1;
   25317: out<=1;
   25318: out<=0;
   25319: out<=0;
   25320: out<=0;
   25321: out<=0;
   25322: out<=0;
   25323: out<=0;
   25324: out<=1;
   25325: out<=0;
   25326: out<=0;
   25327: out<=1;
   25328: out<=0;
   25329: out<=0;
   25330: out<=1;
   25331: out<=1;
   25332: out<=0;
   25333: out<=1;
   25334: out<=0;
   25335: out<=1;
   25336: out<=1;
   25337: out<=0;
   25338: out<=0;
   25339: out<=1;
   25340: out<=1;
   25341: out<=1;
   25342: out<=1;
   25343: out<=1;
   25344: out<=1;
   25345: out<=0;
   25346: out<=0;
   25347: out<=1;
   25348: out<=0;
   25349: out<=0;
   25350: out<=0;
   25351: out<=0;
   25352: out<=0;
   25353: out<=0;
   25354: out<=1;
   25355: out<=1;
   25356: out<=1;
   25357: out<=0;
   25358: out<=1;
   25359: out<=0;
   25360: out<=0;
   25361: out<=0;
   25362: out<=0;
   25363: out<=0;
   25364: out<=0;
   25365: out<=1;
   25366: out<=1;
   25367: out<=0;
   25368: out<=0;
   25369: out<=1;
   25370: out<=0;
   25371: out<=1;
   25372: out<=0;
   25373: out<=0;
   25374: out<=1;
   25375: out<=1;
   25376: out<=0;
   25377: out<=0;
   25378: out<=1;
   25379: out<=1;
   25380: out<=0;
   25381: out<=1;
   25382: out<=0;
   25383: out<=1;
   25384: out<=1;
   25385: out<=0;
   25386: out<=0;
   25387: out<=1;
   25388: out<=1;
   25389: out<=1;
   25390: out<=1;
   25391: out<=1;
   25392: out<=1;
   25393: out<=0;
   25394: out<=1;
   25395: out<=0;
   25396: out<=0;
   25397: out<=0;
   25398: out<=1;
   25399: out<=1;
   25400: out<=1;
   25401: out<=1;
   25402: out<=1;
   25403: out<=1;
   25404: out<=0;
   25405: out<=1;
   25406: out<=1;
   25407: out<=0;
   25408: out<=1;
   25409: out<=0;
   25410: out<=0;
   25411: out<=1;
   25412: out<=0;
   25413: out<=0;
   25414: out<=0;
   25415: out<=0;
   25416: out<=0;
   25417: out<=0;
   25418: out<=1;
   25419: out<=1;
   25420: out<=1;
   25421: out<=0;
   25422: out<=1;
   25423: out<=0;
   25424: out<=1;
   25425: out<=1;
   25426: out<=1;
   25427: out<=1;
   25428: out<=1;
   25429: out<=0;
   25430: out<=0;
   25431: out<=1;
   25432: out<=1;
   25433: out<=0;
   25434: out<=1;
   25435: out<=0;
   25436: out<=1;
   25437: out<=1;
   25438: out<=0;
   25439: out<=0;
   25440: out<=1;
   25441: out<=1;
   25442: out<=0;
   25443: out<=0;
   25444: out<=1;
   25445: out<=0;
   25446: out<=1;
   25447: out<=0;
   25448: out<=0;
   25449: out<=1;
   25450: out<=1;
   25451: out<=0;
   25452: out<=0;
   25453: out<=0;
   25454: out<=0;
   25455: out<=0;
   25456: out<=1;
   25457: out<=0;
   25458: out<=1;
   25459: out<=0;
   25460: out<=0;
   25461: out<=0;
   25462: out<=1;
   25463: out<=1;
   25464: out<=1;
   25465: out<=1;
   25466: out<=1;
   25467: out<=1;
   25468: out<=0;
   25469: out<=1;
   25470: out<=1;
   25471: out<=0;
   25472: out<=1;
   25473: out<=0;
   25474: out<=0;
   25475: out<=1;
   25476: out<=0;
   25477: out<=0;
   25478: out<=0;
   25479: out<=0;
   25480: out<=0;
   25481: out<=0;
   25482: out<=1;
   25483: out<=1;
   25484: out<=1;
   25485: out<=0;
   25486: out<=1;
   25487: out<=0;
   25488: out<=1;
   25489: out<=1;
   25490: out<=1;
   25491: out<=1;
   25492: out<=1;
   25493: out<=0;
   25494: out<=0;
   25495: out<=1;
   25496: out<=1;
   25497: out<=0;
   25498: out<=1;
   25499: out<=0;
   25500: out<=1;
   25501: out<=1;
   25502: out<=0;
   25503: out<=0;
   25504: out<=0;
   25505: out<=0;
   25506: out<=1;
   25507: out<=1;
   25508: out<=0;
   25509: out<=1;
   25510: out<=0;
   25511: out<=1;
   25512: out<=1;
   25513: out<=0;
   25514: out<=0;
   25515: out<=1;
   25516: out<=1;
   25517: out<=1;
   25518: out<=1;
   25519: out<=1;
   25520: out<=0;
   25521: out<=1;
   25522: out<=0;
   25523: out<=1;
   25524: out<=1;
   25525: out<=1;
   25526: out<=0;
   25527: out<=0;
   25528: out<=0;
   25529: out<=0;
   25530: out<=0;
   25531: out<=0;
   25532: out<=1;
   25533: out<=0;
   25534: out<=0;
   25535: out<=1;
   25536: out<=1;
   25537: out<=0;
   25538: out<=0;
   25539: out<=1;
   25540: out<=0;
   25541: out<=0;
   25542: out<=0;
   25543: out<=0;
   25544: out<=0;
   25545: out<=0;
   25546: out<=1;
   25547: out<=1;
   25548: out<=1;
   25549: out<=0;
   25550: out<=1;
   25551: out<=0;
   25552: out<=0;
   25553: out<=0;
   25554: out<=0;
   25555: out<=0;
   25556: out<=0;
   25557: out<=1;
   25558: out<=1;
   25559: out<=0;
   25560: out<=0;
   25561: out<=1;
   25562: out<=0;
   25563: out<=1;
   25564: out<=0;
   25565: out<=0;
   25566: out<=1;
   25567: out<=1;
   25568: out<=1;
   25569: out<=1;
   25570: out<=0;
   25571: out<=0;
   25572: out<=1;
   25573: out<=0;
   25574: out<=1;
   25575: out<=0;
   25576: out<=0;
   25577: out<=1;
   25578: out<=1;
   25579: out<=0;
   25580: out<=0;
   25581: out<=0;
   25582: out<=0;
   25583: out<=0;
   25584: out<=0;
   25585: out<=1;
   25586: out<=0;
   25587: out<=1;
   25588: out<=1;
   25589: out<=1;
   25590: out<=0;
   25591: out<=0;
   25592: out<=0;
   25593: out<=0;
   25594: out<=0;
   25595: out<=0;
   25596: out<=1;
   25597: out<=0;
   25598: out<=0;
   25599: out<=1;
   25600: out<=0;
   25601: out<=0;
   25602: out<=1;
   25603: out<=1;
   25604: out<=1;
   25605: out<=0;
   25606: out<=1;
   25607: out<=0;
   25608: out<=0;
   25609: out<=1;
   25610: out<=1;
   25611: out<=0;
   25612: out<=1;
   25613: out<=1;
   25614: out<=1;
   25615: out<=1;
   25616: out<=1;
   25617: out<=0;
   25618: out<=1;
   25619: out<=0;
   25620: out<=1;
   25621: out<=1;
   25622: out<=0;
   25623: out<=0;
   25624: out<=0;
   25625: out<=0;
   25626: out<=0;
   25627: out<=0;
   25628: out<=0;
   25629: out<=1;
   25630: out<=1;
   25631: out<=0;
   25632: out<=0;
   25633: out<=1;
   25634: out<=1;
   25635: out<=0;
   25636: out<=0;
   25637: out<=0;
   25638: out<=0;
   25639: out<=0;
   25640: out<=0;
   25641: out<=0;
   25642: out<=1;
   25643: out<=1;
   25644: out<=0;
   25645: out<=1;
   25646: out<=0;
   25647: out<=1;
   25648: out<=1;
   25649: out<=1;
   25650: out<=1;
   25651: out<=1;
   25652: out<=0;
   25653: out<=1;
   25654: out<=1;
   25655: out<=0;
   25656: out<=0;
   25657: out<=1;
   25658: out<=0;
   25659: out<=1;
   25660: out<=1;
   25661: out<=1;
   25662: out<=0;
   25663: out<=0;
   25664: out<=1;
   25665: out<=1;
   25666: out<=0;
   25667: out<=0;
   25668: out<=0;
   25669: out<=1;
   25670: out<=0;
   25671: out<=1;
   25672: out<=1;
   25673: out<=0;
   25674: out<=0;
   25675: out<=1;
   25676: out<=0;
   25677: out<=0;
   25678: out<=0;
   25679: out<=0;
   25680: out<=1;
   25681: out<=0;
   25682: out<=1;
   25683: out<=0;
   25684: out<=1;
   25685: out<=1;
   25686: out<=0;
   25687: out<=0;
   25688: out<=0;
   25689: out<=0;
   25690: out<=0;
   25691: out<=0;
   25692: out<=0;
   25693: out<=1;
   25694: out<=1;
   25695: out<=0;
   25696: out<=0;
   25697: out<=1;
   25698: out<=1;
   25699: out<=0;
   25700: out<=0;
   25701: out<=0;
   25702: out<=0;
   25703: out<=0;
   25704: out<=0;
   25705: out<=0;
   25706: out<=1;
   25707: out<=1;
   25708: out<=0;
   25709: out<=1;
   25710: out<=0;
   25711: out<=1;
   25712: out<=0;
   25713: out<=0;
   25714: out<=0;
   25715: out<=0;
   25716: out<=1;
   25717: out<=0;
   25718: out<=0;
   25719: out<=1;
   25720: out<=1;
   25721: out<=0;
   25722: out<=1;
   25723: out<=0;
   25724: out<=0;
   25725: out<=0;
   25726: out<=1;
   25727: out<=1;
   25728: out<=0;
   25729: out<=0;
   25730: out<=1;
   25731: out<=1;
   25732: out<=1;
   25733: out<=0;
   25734: out<=1;
   25735: out<=0;
   25736: out<=0;
   25737: out<=1;
   25738: out<=1;
   25739: out<=0;
   25740: out<=1;
   25741: out<=1;
   25742: out<=1;
   25743: out<=1;
   25744: out<=0;
   25745: out<=1;
   25746: out<=0;
   25747: out<=1;
   25748: out<=0;
   25749: out<=0;
   25750: out<=1;
   25751: out<=1;
   25752: out<=1;
   25753: out<=1;
   25754: out<=1;
   25755: out<=1;
   25756: out<=1;
   25757: out<=0;
   25758: out<=0;
   25759: out<=1;
   25760: out<=0;
   25761: out<=1;
   25762: out<=1;
   25763: out<=0;
   25764: out<=0;
   25765: out<=0;
   25766: out<=0;
   25767: out<=0;
   25768: out<=0;
   25769: out<=0;
   25770: out<=1;
   25771: out<=1;
   25772: out<=0;
   25773: out<=1;
   25774: out<=0;
   25775: out<=1;
   25776: out<=0;
   25777: out<=0;
   25778: out<=0;
   25779: out<=0;
   25780: out<=1;
   25781: out<=0;
   25782: out<=0;
   25783: out<=1;
   25784: out<=1;
   25785: out<=0;
   25786: out<=1;
   25787: out<=0;
   25788: out<=0;
   25789: out<=0;
   25790: out<=1;
   25791: out<=1;
   25792: out<=1;
   25793: out<=1;
   25794: out<=0;
   25795: out<=0;
   25796: out<=0;
   25797: out<=1;
   25798: out<=0;
   25799: out<=1;
   25800: out<=1;
   25801: out<=0;
   25802: out<=0;
   25803: out<=1;
   25804: out<=0;
   25805: out<=0;
   25806: out<=0;
   25807: out<=0;
   25808: out<=0;
   25809: out<=1;
   25810: out<=0;
   25811: out<=1;
   25812: out<=0;
   25813: out<=0;
   25814: out<=1;
   25815: out<=1;
   25816: out<=1;
   25817: out<=1;
   25818: out<=1;
   25819: out<=1;
   25820: out<=1;
   25821: out<=0;
   25822: out<=0;
   25823: out<=1;
   25824: out<=0;
   25825: out<=1;
   25826: out<=1;
   25827: out<=0;
   25828: out<=0;
   25829: out<=0;
   25830: out<=0;
   25831: out<=0;
   25832: out<=0;
   25833: out<=0;
   25834: out<=1;
   25835: out<=1;
   25836: out<=0;
   25837: out<=1;
   25838: out<=0;
   25839: out<=1;
   25840: out<=1;
   25841: out<=1;
   25842: out<=1;
   25843: out<=1;
   25844: out<=0;
   25845: out<=1;
   25846: out<=1;
   25847: out<=0;
   25848: out<=0;
   25849: out<=1;
   25850: out<=0;
   25851: out<=1;
   25852: out<=1;
   25853: out<=1;
   25854: out<=0;
   25855: out<=0;
   25856: out<=1;
   25857: out<=0;
   25858: out<=1;
   25859: out<=0;
   25860: out<=1;
   25861: out<=1;
   25862: out<=0;
   25863: out<=0;
   25864: out<=0;
   25865: out<=0;
   25866: out<=0;
   25867: out<=0;
   25868: out<=0;
   25869: out<=1;
   25870: out<=1;
   25871: out<=0;
   25872: out<=1;
   25873: out<=1;
   25874: out<=0;
   25875: out<=0;
   25876: out<=0;
   25877: out<=1;
   25878: out<=0;
   25879: out<=1;
   25880: out<=1;
   25881: out<=0;
   25882: out<=0;
   25883: out<=1;
   25884: out<=0;
   25885: out<=0;
   25886: out<=0;
   25887: out<=0;
   25888: out<=0;
   25889: out<=0;
   25890: out<=0;
   25891: out<=0;
   25892: out<=1;
   25893: out<=0;
   25894: out<=0;
   25895: out<=1;
   25896: out<=1;
   25897: out<=0;
   25898: out<=1;
   25899: out<=0;
   25900: out<=0;
   25901: out<=0;
   25902: out<=1;
   25903: out<=1;
   25904: out<=0;
   25905: out<=1;
   25906: out<=1;
   25907: out<=0;
   25908: out<=0;
   25909: out<=0;
   25910: out<=0;
   25911: out<=0;
   25912: out<=0;
   25913: out<=0;
   25914: out<=1;
   25915: out<=1;
   25916: out<=0;
   25917: out<=1;
   25918: out<=0;
   25919: out<=1;
   25920: out<=1;
   25921: out<=0;
   25922: out<=1;
   25923: out<=0;
   25924: out<=1;
   25925: out<=1;
   25926: out<=0;
   25927: out<=0;
   25928: out<=0;
   25929: out<=0;
   25930: out<=0;
   25931: out<=0;
   25932: out<=0;
   25933: out<=1;
   25934: out<=1;
   25935: out<=0;
   25936: out<=0;
   25937: out<=0;
   25938: out<=1;
   25939: out<=1;
   25940: out<=1;
   25941: out<=0;
   25942: out<=1;
   25943: out<=0;
   25944: out<=0;
   25945: out<=1;
   25946: out<=1;
   25947: out<=0;
   25948: out<=1;
   25949: out<=1;
   25950: out<=1;
   25951: out<=1;
   25952: out<=1;
   25953: out<=1;
   25954: out<=1;
   25955: out<=1;
   25956: out<=0;
   25957: out<=1;
   25958: out<=1;
   25959: out<=0;
   25960: out<=0;
   25961: out<=1;
   25962: out<=0;
   25963: out<=1;
   25964: out<=1;
   25965: out<=1;
   25966: out<=0;
   25967: out<=0;
   25968: out<=0;
   25969: out<=1;
   25970: out<=1;
   25971: out<=0;
   25972: out<=0;
   25973: out<=0;
   25974: out<=0;
   25975: out<=0;
   25976: out<=0;
   25977: out<=0;
   25978: out<=1;
   25979: out<=1;
   25980: out<=0;
   25981: out<=1;
   25982: out<=0;
   25983: out<=1;
   25984: out<=0;
   25985: out<=1;
   25986: out<=0;
   25987: out<=1;
   25988: out<=0;
   25989: out<=0;
   25990: out<=1;
   25991: out<=1;
   25992: out<=1;
   25993: out<=1;
   25994: out<=1;
   25995: out<=1;
   25996: out<=1;
   25997: out<=0;
   25998: out<=0;
   25999: out<=1;
   26000: out<=1;
   26001: out<=1;
   26002: out<=0;
   26003: out<=0;
   26004: out<=0;
   26005: out<=1;
   26006: out<=0;
   26007: out<=1;
   26008: out<=1;
   26009: out<=0;
   26010: out<=0;
   26011: out<=1;
   26012: out<=0;
   26013: out<=0;
   26014: out<=0;
   26015: out<=0;
   26016: out<=1;
   26017: out<=1;
   26018: out<=1;
   26019: out<=1;
   26020: out<=0;
   26021: out<=1;
   26022: out<=1;
   26023: out<=0;
   26024: out<=0;
   26025: out<=1;
   26026: out<=0;
   26027: out<=1;
   26028: out<=1;
   26029: out<=1;
   26030: out<=0;
   26031: out<=0;
   26032: out<=0;
   26033: out<=1;
   26034: out<=1;
   26035: out<=0;
   26036: out<=0;
   26037: out<=0;
   26038: out<=0;
   26039: out<=0;
   26040: out<=0;
   26041: out<=0;
   26042: out<=1;
   26043: out<=1;
   26044: out<=0;
   26045: out<=1;
   26046: out<=0;
   26047: out<=1;
   26048: out<=0;
   26049: out<=1;
   26050: out<=0;
   26051: out<=1;
   26052: out<=0;
   26053: out<=0;
   26054: out<=1;
   26055: out<=1;
   26056: out<=1;
   26057: out<=1;
   26058: out<=1;
   26059: out<=1;
   26060: out<=1;
   26061: out<=0;
   26062: out<=0;
   26063: out<=1;
   26064: out<=0;
   26065: out<=0;
   26066: out<=1;
   26067: out<=1;
   26068: out<=1;
   26069: out<=0;
   26070: out<=1;
   26071: out<=0;
   26072: out<=0;
   26073: out<=1;
   26074: out<=1;
   26075: out<=0;
   26076: out<=1;
   26077: out<=1;
   26078: out<=1;
   26079: out<=1;
   26080: out<=0;
   26081: out<=0;
   26082: out<=0;
   26083: out<=0;
   26084: out<=1;
   26085: out<=0;
   26086: out<=0;
   26087: out<=1;
   26088: out<=1;
   26089: out<=0;
   26090: out<=1;
   26091: out<=0;
   26092: out<=0;
   26093: out<=0;
   26094: out<=1;
   26095: out<=1;
   26096: out<=0;
   26097: out<=1;
   26098: out<=1;
   26099: out<=0;
   26100: out<=0;
   26101: out<=0;
   26102: out<=0;
   26103: out<=0;
   26104: out<=0;
   26105: out<=0;
   26106: out<=1;
   26107: out<=1;
   26108: out<=0;
   26109: out<=1;
   26110: out<=0;
   26111: out<=1;
   26112: out<=0;
   26113: out<=1;
   26114: out<=1;
   26115: out<=0;
   26116: out<=0;
   26117: out<=0;
   26118: out<=0;
   26119: out<=0;
   26120: out<=0;
   26121: out<=0;
   26122: out<=1;
   26123: out<=1;
   26124: out<=0;
   26125: out<=1;
   26126: out<=0;
   26127: out<=1;
   26128: out<=0;
   26129: out<=0;
   26130: out<=0;
   26131: out<=0;
   26132: out<=1;
   26133: out<=0;
   26134: out<=0;
   26135: out<=1;
   26136: out<=1;
   26137: out<=0;
   26138: out<=1;
   26139: out<=0;
   26140: out<=0;
   26141: out<=0;
   26142: out<=1;
   26143: out<=1;
   26144: out<=0;
   26145: out<=0;
   26146: out<=1;
   26147: out<=1;
   26148: out<=1;
   26149: out<=0;
   26150: out<=1;
   26151: out<=0;
   26152: out<=0;
   26153: out<=1;
   26154: out<=1;
   26155: out<=0;
   26156: out<=1;
   26157: out<=1;
   26158: out<=1;
   26159: out<=1;
   26160: out<=0;
   26161: out<=1;
   26162: out<=0;
   26163: out<=1;
   26164: out<=0;
   26165: out<=0;
   26166: out<=1;
   26167: out<=1;
   26168: out<=1;
   26169: out<=1;
   26170: out<=1;
   26171: out<=1;
   26172: out<=1;
   26173: out<=0;
   26174: out<=0;
   26175: out<=1;
   26176: out<=0;
   26177: out<=1;
   26178: out<=1;
   26179: out<=0;
   26180: out<=0;
   26181: out<=0;
   26182: out<=0;
   26183: out<=0;
   26184: out<=0;
   26185: out<=0;
   26186: out<=1;
   26187: out<=1;
   26188: out<=0;
   26189: out<=1;
   26190: out<=0;
   26191: out<=1;
   26192: out<=1;
   26193: out<=1;
   26194: out<=1;
   26195: out<=1;
   26196: out<=0;
   26197: out<=1;
   26198: out<=1;
   26199: out<=0;
   26200: out<=0;
   26201: out<=1;
   26202: out<=0;
   26203: out<=1;
   26204: out<=1;
   26205: out<=1;
   26206: out<=0;
   26207: out<=0;
   26208: out<=1;
   26209: out<=1;
   26210: out<=0;
   26211: out<=0;
   26212: out<=0;
   26213: out<=1;
   26214: out<=0;
   26215: out<=1;
   26216: out<=1;
   26217: out<=0;
   26218: out<=0;
   26219: out<=1;
   26220: out<=0;
   26221: out<=0;
   26222: out<=0;
   26223: out<=0;
   26224: out<=0;
   26225: out<=1;
   26226: out<=0;
   26227: out<=1;
   26228: out<=0;
   26229: out<=0;
   26230: out<=1;
   26231: out<=1;
   26232: out<=1;
   26233: out<=1;
   26234: out<=1;
   26235: out<=1;
   26236: out<=1;
   26237: out<=0;
   26238: out<=0;
   26239: out<=1;
   26240: out<=0;
   26241: out<=1;
   26242: out<=1;
   26243: out<=0;
   26244: out<=0;
   26245: out<=0;
   26246: out<=0;
   26247: out<=0;
   26248: out<=0;
   26249: out<=0;
   26250: out<=1;
   26251: out<=1;
   26252: out<=0;
   26253: out<=1;
   26254: out<=0;
   26255: out<=1;
   26256: out<=1;
   26257: out<=1;
   26258: out<=1;
   26259: out<=1;
   26260: out<=0;
   26261: out<=1;
   26262: out<=1;
   26263: out<=0;
   26264: out<=0;
   26265: out<=1;
   26266: out<=0;
   26267: out<=1;
   26268: out<=1;
   26269: out<=1;
   26270: out<=0;
   26271: out<=0;
   26272: out<=0;
   26273: out<=0;
   26274: out<=1;
   26275: out<=1;
   26276: out<=1;
   26277: out<=0;
   26278: out<=1;
   26279: out<=0;
   26280: out<=0;
   26281: out<=1;
   26282: out<=1;
   26283: out<=0;
   26284: out<=1;
   26285: out<=1;
   26286: out<=1;
   26287: out<=1;
   26288: out<=1;
   26289: out<=0;
   26290: out<=1;
   26291: out<=0;
   26292: out<=1;
   26293: out<=1;
   26294: out<=0;
   26295: out<=0;
   26296: out<=0;
   26297: out<=0;
   26298: out<=0;
   26299: out<=0;
   26300: out<=0;
   26301: out<=1;
   26302: out<=1;
   26303: out<=0;
   26304: out<=0;
   26305: out<=1;
   26306: out<=1;
   26307: out<=0;
   26308: out<=0;
   26309: out<=0;
   26310: out<=0;
   26311: out<=0;
   26312: out<=0;
   26313: out<=0;
   26314: out<=1;
   26315: out<=1;
   26316: out<=0;
   26317: out<=1;
   26318: out<=0;
   26319: out<=1;
   26320: out<=0;
   26321: out<=0;
   26322: out<=0;
   26323: out<=0;
   26324: out<=1;
   26325: out<=0;
   26326: out<=0;
   26327: out<=1;
   26328: out<=1;
   26329: out<=0;
   26330: out<=1;
   26331: out<=0;
   26332: out<=0;
   26333: out<=0;
   26334: out<=1;
   26335: out<=1;
   26336: out<=1;
   26337: out<=1;
   26338: out<=0;
   26339: out<=0;
   26340: out<=0;
   26341: out<=1;
   26342: out<=0;
   26343: out<=1;
   26344: out<=1;
   26345: out<=0;
   26346: out<=0;
   26347: out<=1;
   26348: out<=0;
   26349: out<=0;
   26350: out<=0;
   26351: out<=0;
   26352: out<=1;
   26353: out<=0;
   26354: out<=1;
   26355: out<=0;
   26356: out<=1;
   26357: out<=1;
   26358: out<=0;
   26359: out<=0;
   26360: out<=0;
   26361: out<=0;
   26362: out<=0;
   26363: out<=0;
   26364: out<=0;
   26365: out<=1;
   26366: out<=1;
   26367: out<=0;
   26368: out<=1;
   26369: out<=1;
   26370: out<=1;
   26371: out<=1;
   26372: out<=0;
   26373: out<=1;
   26374: out<=1;
   26375: out<=0;
   26376: out<=0;
   26377: out<=1;
   26378: out<=0;
   26379: out<=1;
   26380: out<=1;
   26381: out<=1;
   26382: out<=0;
   26383: out<=0;
   26384: out<=0;
   26385: out<=1;
   26386: out<=1;
   26387: out<=0;
   26388: out<=0;
   26389: out<=0;
   26390: out<=0;
   26391: out<=0;
   26392: out<=0;
   26393: out<=0;
   26394: out<=1;
   26395: out<=1;
   26396: out<=0;
   26397: out<=1;
   26398: out<=0;
   26399: out<=1;
   26400: out<=0;
   26401: out<=1;
   26402: out<=0;
   26403: out<=1;
   26404: out<=0;
   26405: out<=0;
   26406: out<=1;
   26407: out<=1;
   26408: out<=1;
   26409: out<=1;
   26410: out<=1;
   26411: out<=1;
   26412: out<=1;
   26413: out<=0;
   26414: out<=0;
   26415: out<=1;
   26416: out<=1;
   26417: out<=1;
   26418: out<=0;
   26419: out<=0;
   26420: out<=0;
   26421: out<=1;
   26422: out<=0;
   26423: out<=1;
   26424: out<=1;
   26425: out<=0;
   26426: out<=0;
   26427: out<=1;
   26428: out<=0;
   26429: out<=0;
   26430: out<=0;
   26431: out<=0;
   26432: out<=0;
   26433: out<=0;
   26434: out<=0;
   26435: out<=0;
   26436: out<=1;
   26437: out<=0;
   26438: out<=0;
   26439: out<=1;
   26440: out<=1;
   26441: out<=0;
   26442: out<=1;
   26443: out<=0;
   26444: out<=0;
   26445: out<=0;
   26446: out<=1;
   26447: out<=1;
   26448: out<=0;
   26449: out<=1;
   26450: out<=1;
   26451: out<=0;
   26452: out<=0;
   26453: out<=0;
   26454: out<=0;
   26455: out<=0;
   26456: out<=0;
   26457: out<=0;
   26458: out<=1;
   26459: out<=1;
   26460: out<=0;
   26461: out<=1;
   26462: out<=0;
   26463: out<=1;
   26464: out<=0;
   26465: out<=1;
   26466: out<=0;
   26467: out<=1;
   26468: out<=0;
   26469: out<=0;
   26470: out<=1;
   26471: out<=1;
   26472: out<=1;
   26473: out<=1;
   26474: out<=1;
   26475: out<=1;
   26476: out<=1;
   26477: out<=0;
   26478: out<=0;
   26479: out<=1;
   26480: out<=0;
   26481: out<=0;
   26482: out<=1;
   26483: out<=1;
   26484: out<=1;
   26485: out<=0;
   26486: out<=1;
   26487: out<=0;
   26488: out<=0;
   26489: out<=1;
   26490: out<=1;
   26491: out<=0;
   26492: out<=1;
   26493: out<=1;
   26494: out<=1;
   26495: out<=1;
   26496: out<=0;
   26497: out<=0;
   26498: out<=0;
   26499: out<=0;
   26500: out<=1;
   26501: out<=0;
   26502: out<=0;
   26503: out<=1;
   26504: out<=1;
   26505: out<=0;
   26506: out<=1;
   26507: out<=0;
   26508: out<=0;
   26509: out<=0;
   26510: out<=1;
   26511: out<=1;
   26512: out<=0;
   26513: out<=1;
   26514: out<=1;
   26515: out<=0;
   26516: out<=0;
   26517: out<=0;
   26518: out<=0;
   26519: out<=0;
   26520: out<=0;
   26521: out<=0;
   26522: out<=1;
   26523: out<=1;
   26524: out<=0;
   26525: out<=1;
   26526: out<=0;
   26527: out<=1;
   26528: out<=1;
   26529: out<=0;
   26530: out<=1;
   26531: out<=0;
   26532: out<=1;
   26533: out<=1;
   26534: out<=0;
   26535: out<=0;
   26536: out<=0;
   26537: out<=0;
   26538: out<=0;
   26539: out<=0;
   26540: out<=0;
   26541: out<=1;
   26542: out<=1;
   26543: out<=0;
   26544: out<=1;
   26545: out<=1;
   26546: out<=0;
   26547: out<=0;
   26548: out<=0;
   26549: out<=1;
   26550: out<=0;
   26551: out<=1;
   26552: out<=1;
   26553: out<=0;
   26554: out<=0;
   26555: out<=1;
   26556: out<=0;
   26557: out<=0;
   26558: out<=0;
   26559: out<=0;
   26560: out<=1;
   26561: out<=1;
   26562: out<=1;
   26563: out<=1;
   26564: out<=0;
   26565: out<=1;
   26566: out<=1;
   26567: out<=0;
   26568: out<=0;
   26569: out<=1;
   26570: out<=0;
   26571: out<=1;
   26572: out<=1;
   26573: out<=1;
   26574: out<=0;
   26575: out<=0;
   26576: out<=0;
   26577: out<=1;
   26578: out<=1;
   26579: out<=0;
   26580: out<=0;
   26581: out<=0;
   26582: out<=0;
   26583: out<=0;
   26584: out<=0;
   26585: out<=0;
   26586: out<=1;
   26587: out<=1;
   26588: out<=0;
   26589: out<=1;
   26590: out<=0;
   26591: out<=1;
   26592: out<=1;
   26593: out<=0;
   26594: out<=1;
   26595: out<=0;
   26596: out<=1;
   26597: out<=1;
   26598: out<=0;
   26599: out<=0;
   26600: out<=0;
   26601: out<=0;
   26602: out<=0;
   26603: out<=0;
   26604: out<=0;
   26605: out<=1;
   26606: out<=1;
   26607: out<=0;
   26608: out<=0;
   26609: out<=0;
   26610: out<=1;
   26611: out<=1;
   26612: out<=1;
   26613: out<=0;
   26614: out<=1;
   26615: out<=0;
   26616: out<=0;
   26617: out<=1;
   26618: out<=1;
   26619: out<=0;
   26620: out<=1;
   26621: out<=1;
   26622: out<=1;
   26623: out<=1;
   26624: out<=1;
   26625: out<=1;
   26626: out<=1;
   26627: out<=1;
   26628: out<=0;
   26629: out<=1;
   26630: out<=1;
   26631: out<=0;
   26632: out<=1;
   26633: out<=0;
   26634: out<=1;
   26635: out<=0;
   26636: out<=0;
   26637: out<=0;
   26638: out<=1;
   26639: out<=1;
   26640: out<=0;
   26641: out<=1;
   26642: out<=1;
   26643: out<=0;
   26644: out<=0;
   26645: out<=0;
   26646: out<=0;
   26647: out<=0;
   26648: out<=1;
   26649: out<=1;
   26650: out<=0;
   26651: out<=0;
   26652: out<=1;
   26653: out<=0;
   26654: out<=1;
   26655: out<=0;
   26656: out<=1;
   26657: out<=0;
   26658: out<=1;
   26659: out<=0;
   26660: out<=1;
   26661: out<=1;
   26662: out<=0;
   26663: out<=0;
   26664: out<=1;
   26665: out<=1;
   26666: out<=1;
   26667: out<=1;
   26668: out<=1;
   26669: out<=0;
   26670: out<=0;
   26671: out<=1;
   26672: out<=0;
   26673: out<=0;
   26674: out<=1;
   26675: out<=1;
   26676: out<=1;
   26677: out<=0;
   26678: out<=1;
   26679: out<=0;
   26680: out<=1;
   26681: out<=0;
   26682: out<=0;
   26683: out<=1;
   26684: out<=0;
   26685: out<=0;
   26686: out<=0;
   26687: out<=0;
   26688: out<=0;
   26689: out<=0;
   26690: out<=0;
   26691: out<=0;
   26692: out<=1;
   26693: out<=0;
   26694: out<=0;
   26695: out<=1;
   26696: out<=0;
   26697: out<=1;
   26698: out<=0;
   26699: out<=1;
   26700: out<=1;
   26701: out<=1;
   26702: out<=0;
   26703: out<=0;
   26704: out<=0;
   26705: out<=1;
   26706: out<=1;
   26707: out<=0;
   26708: out<=0;
   26709: out<=0;
   26710: out<=0;
   26711: out<=0;
   26712: out<=1;
   26713: out<=1;
   26714: out<=0;
   26715: out<=0;
   26716: out<=1;
   26717: out<=0;
   26718: out<=1;
   26719: out<=0;
   26720: out<=1;
   26721: out<=0;
   26722: out<=1;
   26723: out<=0;
   26724: out<=1;
   26725: out<=1;
   26726: out<=0;
   26727: out<=0;
   26728: out<=1;
   26729: out<=1;
   26730: out<=1;
   26731: out<=1;
   26732: out<=1;
   26733: out<=0;
   26734: out<=0;
   26735: out<=1;
   26736: out<=1;
   26737: out<=1;
   26738: out<=0;
   26739: out<=0;
   26740: out<=0;
   26741: out<=1;
   26742: out<=0;
   26743: out<=1;
   26744: out<=0;
   26745: out<=1;
   26746: out<=1;
   26747: out<=0;
   26748: out<=1;
   26749: out<=1;
   26750: out<=1;
   26751: out<=1;
   26752: out<=0;
   26753: out<=0;
   26754: out<=0;
   26755: out<=0;
   26756: out<=1;
   26757: out<=0;
   26758: out<=0;
   26759: out<=1;
   26760: out<=0;
   26761: out<=1;
   26762: out<=0;
   26763: out<=1;
   26764: out<=1;
   26765: out<=1;
   26766: out<=0;
   26767: out<=0;
   26768: out<=0;
   26769: out<=1;
   26770: out<=1;
   26771: out<=0;
   26772: out<=0;
   26773: out<=0;
   26774: out<=0;
   26775: out<=0;
   26776: out<=1;
   26777: out<=1;
   26778: out<=0;
   26779: out<=0;
   26780: out<=1;
   26781: out<=0;
   26782: out<=1;
   26783: out<=0;
   26784: out<=0;
   26785: out<=1;
   26786: out<=0;
   26787: out<=1;
   26788: out<=0;
   26789: out<=0;
   26790: out<=1;
   26791: out<=1;
   26792: out<=0;
   26793: out<=0;
   26794: out<=0;
   26795: out<=0;
   26796: out<=0;
   26797: out<=1;
   26798: out<=1;
   26799: out<=0;
   26800: out<=0;
   26801: out<=0;
   26802: out<=1;
   26803: out<=1;
   26804: out<=1;
   26805: out<=0;
   26806: out<=1;
   26807: out<=0;
   26808: out<=1;
   26809: out<=0;
   26810: out<=0;
   26811: out<=1;
   26812: out<=0;
   26813: out<=0;
   26814: out<=0;
   26815: out<=0;
   26816: out<=1;
   26817: out<=1;
   26818: out<=1;
   26819: out<=1;
   26820: out<=0;
   26821: out<=1;
   26822: out<=1;
   26823: out<=0;
   26824: out<=1;
   26825: out<=0;
   26826: out<=1;
   26827: out<=0;
   26828: out<=0;
   26829: out<=0;
   26830: out<=1;
   26831: out<=1;
   26832: out<=0;
   26833: out<=1;
   26834: out<=1;
   26835: out<=0;
   26836: out<=0;
   26837: out<=0;
   26838: out<=0;
   26839: out<=0;
   26840: out<=1;
   26841: out<=1;
   26842: out<=0;
   26843: out<=0;
   26844: out<=1;
   26845: out<=0;
   26846: out<=1;
   26847: out<=0;
   26848: out<=0;
   26849: out<=1;
   26850: out<=0;
   26851: out<=1;
   26852: out<=0;
   26853: out<=0;
   26854: out<=1;
   26855: out<=1;
   26856: out<=0;
   26857: out<=0;
   26858: out<=0;
   26859: out<=0;
   26860: out<=0;
   26861: out<=1;
   26862: out<=1;
   26863: out<=0;
   26864: out<=1;
   26865: out<=1;
   26866: out<=0;
   26867: out<=0;
   26868: out<=0;
   26869: out<=1;
   26870: out<=0;
   26871: out<=1;
   26872: out<=0;
   26873: out<=1;
   26874: out<=1;
   26875: out<=0;
   26876: out<=1;
   26877: out<=1;
   26878: out<=1;
   26879: out<=1;
   26880: out<=0;
   26881: out<=1;
   26882: out<=1;
   26883: out<=0;
   26884: out<=0;
   26885: out<=0;
   26886: out<=0;
   26887: out<=0;
   26888: out<=1;
   26889: out<=1;
   26890: out<=0;
   26891: out<=0;
   26892: out<=1;
   26893: out<=0;
   26894: out<=1;
   26895: out<=0;
   26896: out<=0;
   26897: out<=0;
   26898: out<=0;
   26899: out<=0;
   26900: out<=1;
   26901: out<=0;
   26902: out<=0;
   26903: out<=1;
   26904: out<=0;
   26905: out<=1;
   26906: out<=0;
   26907: out<=1;
   26908: out<=1;
   26909: out<=1;
   26910: out<=0;
   26911: out<=0;
   26912: out<=1;
   26913: out<=1;
   26914: out<=0;
   26915: out<=0;
   26916: out<=0;
   26917: out<=1;
   26918: out<=0;
   26919: out<=1;
   26920: out<=0;
   26921: out<=1;
   26922: out<=1;
   26923: out<=0;
   26924: out<=1;
   26925: out<=1;
   26926: out<=1;
   26927: out<=1;
   26928: out<=1;
   26929: out<=0;
   26930: out<=1;
   26931: out<=0;
   26932: out<=1;
   26933: out<=1;
   26934: out<=0;
   26935: out<=0;
   26936: out<=1;
   26937: out<=1;
   26938: out<=1;
   26939: out<=1;
   26940: out<=1;
   26941: out<=0;
   26942: out<=0;
   26943: out<=1;
   26944: out<=0;
   26945: out<=1;
   26946: out<=1;
   26947: out<=0;
   26948: out<=0;
   26949: out<=0;
   26950: out<=0;
   26951: out<=0;
   26952: out<=1;
   26953: out<=1;
   26954: out<=0;
   26955: out<=0;
   26956: out<=1;
   26957: out<=0;
   26958: out<=1;
   26959: out<=0;
   26960: out<=1;
   26961: out<=1;
   26962: out<=1;
   26963: out<=1;
   26964: out<=0;
   26965: out<=1;
   26966: out<=1;
   26967: out<=0;
   26968: out<=1;
   26969: out<=0;
   26970: out<=1;
   26971: out<=0;
   26972: out<=0;
   26973: out<=0;
   26974: out<=1;
   26975: out<=1;
   26976: out<=0;
   26977: out<=0;
   26978: out<=1;
   26979: out<=1;
   26980: out<=1;
   26981: out<=0;
   26982: out<=1;
   26983: out<=0;
   26984: out<=1;
   26985: out<=0;
   26986: out<=0;
   26987: out<=1;
   26988: out<=0;
   26989: out<=0;
   26990: out<=0;
   26991: out<=0;
   26992: out<=1;
   26993: out<=0;
   26994: out<=1;
   26995: out<=0;
   26996: out<=1;
   26997: out<=1;
   26998: out<=0;
   26999: out<=0;
   27000: out<=1;
   27001: out<=1;
   27002: out<=1;
   27003: out<=1;
   27004: out<=1;
   27005: out<=0;
   27006: out<=0;
   27007: out<=1;
   27008: out<=0;
   27009: out<=1;
   27010: out<=1;
   27011: out<=0;
   27012: out<=0;
   27013: out<=0;
   27014: out<=0;
   27015: out<=0;
   27016: out<=1;
   27017: out<=1;
   27018: out<=0;
   27019: out<=0;
   27020: out<=1;
   27021: out<=0;
   27022: out<=1;
   27023: out<=0;
   27024: out<=1;
   27025: out<=1;
   27026: out<=1;
   27027: out<=1;
   27028: out<=0;
   27029: out<=1;
   27030: out<=1;
   27031: out<=0;
   27032: out<=1;
   27033: out<=0;
   27034: out<=1;
   27035: out<=0;
   27036: out<=0;
   27037: out<=0;
   27038: out<=1;
   27039: out<=1;
   27040: out<=1;
   27041: out<=1;
   27042: out<=0;
   27043: out<=0;
   27044: out<=0;
   27045: out<=1;
   27046: out<=0;
   27047: out<=1;
   27048: out<=0;
   27049: out<=1;
   27050: out<=1;
   27051: out<=0;
   27052: out<=1;
   27053: out<=1;
   27054: out<=1;
   27055: out<=1;
   27056: out<=0;
   27057: out<=1;
   27058: out<=0;
   27059: out<=1;
   27060: out<=0;
   27061: out<=0;
   27062: out<=1;
   27063: out<=1;
   27064: out<=0;
   27065: out<=0;
   27066: out<=0;
   27067: out<=0;
   27068: out<=0;
   27069: out<=1;
   27070: out<=1;
   27071: out<=0;
   27072: out<=0;
   27073: out<=1;
   27074: out<=1;
   27075: out<=0;
   27076: out<=0;
   27077: out<=0;
   27078: out<=0;
   27079: out<=0;
   27080: out<=1;
   27081: out<=1;
   27082: out<=0;
   27083: out<=0;
   27084: out<=1;
   27085: out<=0;
   27086: out<=1;
   27087: out<=0;
   27088: out<=0;
   27089: out<=0;
   27090: out<=0;
   27091: out<=0;
   27092: out<=1;
   27093: out<=0;
   27094: out<=0;
   27095: out<=1;
   27096: out<=0;
   27097: out<=1;
   27098: out<=0;
   27099: out<=1;
   27100: out<=1;
   27101: out<=1;
   27102: out<=0;
   27103: out<=0;
   27104: out<=0;
   27105: out<=0;
   27106: out<=1;
   27107: out<=1;
   27108: out<=1;
   27109: out<=0;
   27110: out<=1;
   27111: out<=0;
   27112: out<=1;
   27113: out<=0;
   27114: out<=0;
   27115: out<=1;
   27116: out<=0;
   27117: out<=0;
   27118: out<=0;
   27119: out<=0;
   27120: out<=0;
   27121: out<=1;
   27122: out<=0;
   27123: out<=1;
   27124: out<=0;
   27125: out<=0;
   27126: out<=1;
   27127: out<=1;
   27128: out<=0;
   27129: out<=0;
   27130: out<=0;
   27131: out<=0;
   27132: out<=0;
   27133: out<=1;
   27134: out<=1;
   27135: out<=0;
   27136: out<=0;
   27137: out<=1;
   27138: out<=0;
   27139: out<=1;
   27140: out<=0;
   27141: out<=0;
   27142: out<=1;
   27143: out<=1;
   27144: out<=0;
   27145: out<=0;
   27146: out<=0;
   27147: out<=0;
   27148: out<=0;
   27149: out<=1;
   27150: out<=1;
   27151: out<=0;
   27152: out<=0;
   27153: out<=0;
   27154: out<=1;
   27155: out<=1;
   27156: out<=1;
   27157: out<=0;
   27158: out<=1;
   27159: out<=0;
   27160: out<=1;
   27161: out<=0;
   27162: out<=0;
   27163: out<=1;
   27164: out<=0;
   27165: out<=0;
   27166: out<=0;
   27167: out<=0;
   27168: out<=0;
   27169: out<=0;
   27170: out<=0;
   27171: out<=0;
   27172: out<=1;
   27173: out<=0;
   27174: out<=0;
   27175: out<=1;
   27176: out<=0;
   27177: out<=1;
   27178: out<=0;
   27179: out<=1;
   27180: out<=1;
   27181: out<=1;
   27182: out<=0;
   27183: out<=0;
   27184: out<=0;
   27185: out<=1;
   27186: out<=1;
   27187: out<=0;
   27188: out<=0;
   27189: out<=0;
   27190: out<=0;
   27191: out<=0;
   27192: out<=1;
   27193: out<=1;
   27194: out<=0;
   27195: out<=0;
   27196: out<=1;
   27197: out<=0;
   27198: out<=1;
   27199: out<=0;
   27200: out<=0;
   27201: out<=1;
   27202: out<=0;
   27203: out<=1;
   27204: out<=0;
   27205: out<=0;
   27206: out<=1;
   27207: out<=1;
   27208: out<=0;
   27209: out<=0;
   27210: out<=0;
   27211: out<=0;
   27212: out<=0;
   27213: out<=1;
   27214: out<=1;
   27215: out<=0;
   27216: out<=1;
   27217: out<=1;
   27218: out<=0;
   27219: out<=0;
   27220: out<=0;
   27221: out<=1;
   27222: out<=0;
   27223: out<=1;
   27224: out<=0;
   27225: out<=1;
   27226: out<=1;
   27227: out<=0;
   27228: out<=1;
   27229: out<=1;
   27230: out<=1;
   27231: out<=1;
   27232: out<=1;
   27233: out<=1;
   27234: out<=1;
   27235: out<=1;
   27236: out<=0;
   27237: out<=1;
   27238: out<=1;
   27239: out<=0;
   27240: out<=1;
   27241: out<=0;
   27242: out<=1;
   27243: out<=0;
   27244: out<=0;
   27245: out<=0;
   27246: out<=1;
   27247: out<=1;
   27248: out<=0;
   27249: out<=1;
   27250: out<=1;
   27251: out<=0;
   27252: out<=0;
   27253: out<=0;
   27254: out<=0;
   27255: out<=0;
   27256: out<=1;
   27257: out<=1;
   27258: out<=0;
   27259: out<=0;
   27260: out<=1;
   27261: out<=0;
   27262: out<=1;
   27263: out<=0;
   27264: out<=1;
   27265: out<=0;
   27266: out<=1;
   27267: out<=0;
   27268: out<=1;
   27269: out<=1;
   27270: out<=0;
   27271: out<=0;
   27272: out<=1;
   27273: out<=1;
   27274: out<=1;
   27275: out<=1;
   27276: out<=1;
   27277: out<=0;
   27278: out<=0;
   27279: out<=1;
   27280: out<=0;
   27281: out<=0;
   27282: out<=1;
   27283: out<=1;
   27284: out<=1;
   27285: out<=0;
   27286: out<=1;
   27287: out<=0;
   27288: out<=1;
   27289: out<=0;
   27290: out<=0;
   27291: out<=1;
   27292: out<=0;
   27293: out<=0;
   27294: out<=0;
   27295: out<=0;
   27296: out<=1;
   27297: out<=1;
   27298: out<=1;
   27299: out<=1;
   27300: out<=0;
   27301: out<=1;
   27302: out<=1;
   27303: out<=0;
   27304: out<=1;
   27305: out<=0;
   27306: out<=1;
   27307: out<=0;
   27308: out<=0;
   27309: out<=0;
   27310: out<=1;
   27311: out<=1;
   27312: out<=0;
   27313: out<=1;
   27314: out<=1;
   27315: out<=0;
   27316: out<=0;
   27317: out<=0;
   27318: out<=0;
   27319: out<=0;
   27320: out<=1;
   27321: out<=1;
   27322: out<=0;
   27323: out<=0;
   27324: out<=1;
   27325: out<=0;
   27326: out<=1;
   27327: out<=0;
   27328: out<=1;
   27329: out<=0;
   27330: out<=1;
   27331: out<=0;
   27332: out<=1;
   27333: out<=1;
   27334: out<=0;
   27335: out<=0;
   27336: out<=1;
   27337: out<=1;
   27338: out<=1;
   27339: out<=1;
   27340: out<=1;
   27341: out<=0;
   27342: out<=0;
   27343: out<=1;
   27344: out<=1;
   27345: out<=1;
   27346: out<=0;
   27347: out<=0;
   27348: out<=0;
   27349: out<=1;
   27350: out<=0;
   27351: out<=1;
   27352: out<=0;
   27353: out<=1;
   27354: out<=1;
   27355: out<=0;
   27356: out<=1;
   27357: out<=1;
   27358: out<=1;
   27359: out<=1;
   27360: out<=0;
   27361: out<=0;
   27362: out<=0;
   27363: out<=0;
   27364: out<=1;
   27365: out<=0;
   27366: out<=0;
   27367: out<=1;
   27368: out<=0;
   27369: out<=1;
   27370: out<=0;
   27371: out<=1;
   27372: out<=1;
   27373: out<=1;
   27374: out<=0;
   27375: out<=0;
   27376: out<=0;
   27377: out<=1;
   27378: out<=1;
   27379: out<=0;
   27380: out<=0;
   27381: out<=0;
   27382: out<=0;
   27383: out<=0;
   27384: out<=1;
   27385: out<=1;
   27386: out<=0;
   27387: out<=0;
   27388: out<=1;
   27389: out<=0;
   27390: out<=1;
   27391: out<=0;
   27392: out<=1;
   27393: out<=1;
   27394: out<=0;
   27395: out<=0;
   27396: out<=0;
   27397: out<=1;
   27398: out<=0;
   27399: out<=1;
   27400: out<=0;
   27401: out<=1;
   27402: out<=1;
   27403: out<=0;
   27404: out<=1;
   27405: out<=1;
   27406: out<=1;
   27407: out<=1;
   27408: out<=0;
   27409: out<=1;
   27410: out<=0;
   27411: out<=1;
   27412: out<=0;
   27413: out<=0;
   27414: out<=1;
   27415: out<=1;
   27416: out<=0;
   27417: out<=0;
   27418: out<=0;
   27419: out<=0;
   27420: out<=0;
   27421: out<=1;
   27422: out<=1;
   27423: out<=0;
   27424: out<=0;
   27425: out<=1;
   27426: out<=1;
   27427: out<=0;
   27428: out<=0;
   27429: out<=0;
   27430: out<=0;
   27431: out<=0;
   27432: out<=1;
   27433: out<=1;
   27434: out<=0;
   27435: out<=0;
   27436: out<=1;
   27437: out<=0;
   27438: out<=1;
   27439: out<=0;
   27440: out<=1;
   27441: out<=1;
   27442: out<=1;
   27443: out<=1;
   27444: out<=0;
   27445: out<=1;
   27446: out<=1;
   27447: out<=0;
   27448: out<=1;
   27449: out<=0;
   27450: out<=1;
   27451: out<=0;
   27452: out<=0;
   27453: out<=0;
   27454: out<=1;
   27455: out<=1;
   27456: out<=0;
   27457: out<=0;
   27458: out<=1;
   27459: out<=1;
   27460: out<=1;
   27461: out<=0;
   27462: out<=1;
   27463: out<=0;
   27464: out<=1;
   27465: out<=0;
   27466: out<=0;
   27467: out<=1;
   27468: out<=0;
   27469: out<=0;
   27470: out<=0;
   27471: out<=0;
   27472: out<=0;
   27473: out<=1;
   27474: out<=0;
   27475: out<=1;
   27476: out<=0;
   27477: out<=0;
   27478: out<=1;
   27479: out<=1;
   27480: out<=0;
   27481: out<=0;
   27482: out<=0;
   27483: out<=0;
   27484: out<=0;
   27485: out<=1;
   27486: out<=1;
   27487: out<=0;
   27488: out<=0;
   27489: out<=1;
   27490: out<=1;
   27491: out<=0;
   27492: out<=0;
   27493: out<=0;
   27494: out<=0;
   27495: out<=0;
   27496: out<=1;
   27497: out<=1;
   27498: out<=0;
   27499: out<=0;
   27500: out<=1;
   27501: out<=0;
   27502: out<=1;
   27503: out<=0;
   27504: out<=0;
   27505: out<=0;
   27506: out<=0;
   27507: out<=0;
   27508: out<=1;
   27509: out<=0;
   27510: out<=0;
   27511: out<=1;
   27512: out<=0;
   27513: out<=1;
   27514: out<=0;
   27515: out<=1;
   27516: out<=1;
   27517: out<=1;
   27518: out<=0;
   27519: out<=0;
   27520: out<=1;
   27521: out<=1;
   27522: out<=0;
   27523: out<=0;
   27524: out<=0;
   27525: out<=1;
   27526: out<=0;
   27527: out<=1;
   27528: out<=0;
   27529: out<=1;
   27530: out<=1;
   27531: out<=0;
   27532: out<=1;
   27533: out<=1;
   27534: out<=1;
   27535: out<=1;
   27536: out<=1;
   27537: out<=0;
   27538: out<=1;
   27539: out<=0;
   27540: out<=1;
   27541: out<=1;
   27542: out<=0;
   27543: out<=0;
   27544: out<=1;
   27545: out<=1;
   27546: out<=1;
   27547: out<=1;
   27548: out<=1;
   27549: out<=0;
   27550: out<=0;
   27551: out<=1;
   27552: out<=0;
   27553: out<=1;
   27554: out<=1;
   27555: out<=0;
   27556: out<=0;
   27557: out<=0;
   27558: out<=0;
   27559: out<=0;
   27560: out<=1;
   27561: out<=1;
   27562: out<=0;
   27563: out<=0;
   27564: out<=1;
   27565: out<=0;
   27566: out<=1;
   27567: out<=0;
   27568: out<=0;
   27569: out<=0;
   27570: out<=0;
   27571: out<=0;
   27572: out<=1;
   27573: out<=0;
   27574: out<=0;
   27575: out<=1;
   27576: out<=0;
   27577: out<=1;
   27578: out<=0;
   27579: out<=1;
   27580: out<=1;
   27581: out<=1;
   27582: out<=0;
   27583: out<=0;
   27584: out<=0;
   27585: out<=0;
   27586: out<=1;
   27587: out<=1;
   27588: out<=1;
   27589: out<=0;
   27590: out<=1;
   27591: out<=0;
   27592: out<=1;
   27593: out<=0;
   27594: out<=0;
   27595: out<=1;
   27596: out<=0;
   27597: out<=0;
   27598: out<=0;
   27599: out<=0;
   27600: out<=1;
   27601: out<=0;
   27602: out<=1;
   27603: out<=0;
   27604: out<=1;
   27605: out<=1;
   27606: out<=0;
   27607: out<=0;
   27608: out<=1;
   27609: out<=1;
   27610: out<=1;
   27611: out<=1;
   27612: out<=1;
   27613: out<=0;
   27614: out<=0;
   27615: out<=1;
   27616: out<=0;
   27617: out<=1;
   27618: out<=1;
   27619: out<=0;
   27620: out<=0;
   27621: out<=0;
   27622: out<=0;
   27623: out<=0;
   27624: out<=1;
   27625: out<=1;
   27626: out<=0;
   27627: out<=0;
   27628: out<=1;
   27629: out<=0;
   27630: out<=1;
   27631: out<=0;
   27632: out<=1;
   27633: out<=1;
   27634: out<=1;
   27635: out<=1;
   27636: out<=0;
   27637: out<=1;
   27638: out<=1;
   27639: out<=0;
   27640: out<=1;
   27641: out<=0;
   27642: out<=1;
   27643: out<=0;
   27644: out<=0;
   27645: out<=0;
   27646: out<=1;
   27647: out<=1;
   27648: out<=1;
   27649: out<=0;
   27650: out<=0;
   27651: out<=1;
   27652: out<=0;
   27653: out<=0;
   27654: out<=0;
   27655: out<=0;
   27656: out<=1;
   27657: out<=1;
   27658: out<=0;
   27659: out<=0;
   27660: out<=0;
   27661: out<=1;
   27662: out<=0;
   27663: out<=1;
   27664: out<=0;
   27665: out<=0;
   27666: out<=0;
   27667: out<=0;
   27668: out<=0;
   27669: out<=1;
   27670: out<=1;
   27671: out<=0;
   27672: out<=1;
   27673: out<=0;
   27674: out<=1;
   27675: out<=0;
   27676: out<=1;
   27677: out<=1;
   27678: out<=0;
   27679: out<=0;
   27680: out<=1;
   27681: out<=1;
   27682: out<=0;
   27683: out<=0;
   27684: out<=1;
   27685: out<=0;
   27686: out<=1;
   27687: out<=0;
   27688: out<=1;
   27689: out<=0;
   27690: out<=0;
   27691: out<=1;
   27692: out<=1;
   27693: out<=1;
   27694: out<=1;
   27695: out<=1;
   27696: out<=0;
   27697: out<=1;
   27698: out<=0;
   27699: out<=1;
   27700: out<=1;
   27701: out<=1;
   27702: out<=0;
   27703: out<=0;
   27704: out<=1;
   27705: out<=1;
   27706: out<=1;
   27707: out<=1;
   27708: out<=0;
   27709: out<=1;
   27710: out<=1;
   27711: out<=0;
   27712: out<=1;
   27713: out<=0;
   27714: out<=0;
   27715: out<=1;
   27716: out<=0;
   27717: out<=0;
   27718: out<=0;
   27719: out<=0;
   27720: out<=1;
   27721: out<=1;
   27722: out<=0;
   27723: out<=0;
   27724: out<=0;
   27725: out<=1;
   27726: out<=0;
   27727: out<=1;
   27728: out<=1;
   27729: out<=1;
   27730: out<=1;
   27731: out<=1;
   27732: out<=1;
   27733: out<=0;
   27734: out<=0;
   27735: out<=1;
   27736: out<=0;
   27737: out<=1;
   27738: out<=0;
   27739: out<=1;
   27740: out<=0;
   27741: out<=0;
   27742: out<=1;
   27743: out<=1;
   27744: out<=0;
   27745: out<=0;
   27746: out<=1;
   27747: out<=1;
   27748: out<=0;
   27749: out<=1;
   27750: out<=0;
   27751: out<=1;
   27752: out<=0;
   27753: out<=1;
   27754: out<=1;
   27755: out<=0;
   27756: out<=0;
   27757: out<=0;
   27758: out<=0;
   27759: out<=0;
   27760: out<=0;
   27761: out<=1;
   27762: out<=0;
   27763: out<=1;
   27764: out<=1;
   27765: out<=1;
   27766: out<=0;
   27767: out<=0;
   27768: out<=1;
   27769: out<=1;
   27770: out<=1;
   27771: out<=1;
   27772: out<=0;
   27773: out<=1;
   27774: out<=1;
   27775: out<=0;
   27776: out<=1;
   27777: out<=0;
   27778: out<=0;
   27779: out<=1;
   27780: out<=0;
   27781: out<=0;
   27782: out<=0;
   27783: out<=0;
   27784: out<=1;
   27785: out<=1;
   27786: out<=0;
   27787: out<=0;
   27788: out<=0;
   27789: out<=1;
   27790: out<=0;
   27791: out<=1;
   27792: out<=1;
   27793: out<=1;
   27794: out<=1;
   27795: out<=1;
   27796: out<=1;
   27797: out<=0;
   27798: out<=0;
   27799: out<=1;
   27800: out<=0;
   27801: out<=1;
   27802: out<=0;
   27803: out<=1;
   27804: out<=0;
   27805: out<=0;
   27806: out<=1;
   27807: out<=1;
   27808: out<=1;
   27809: out<=1;
   27810: out<=0;
   27811: out<=0;
   27812: out<=1;
   27813: out<=0;
   27814: out<=1;
   27815: out<=0;
   27816: out<=1;
   27817: out<=0;
   27818: out<=0;
   27819: out<=1;
   27820: out<=1;
   27821: out<=1;
   27822: out<=1;
   27823: out<=1;
   27824: out<=1;
   27825: out<=0;
   27826: out<=1;
   27827: out<=0;
   27828: out<=0;
   27829: out<=0;
   27830: out<=1;
   27831: out<=1;
   27832: out<=0;
   27833: out<=0;
   27834: out<=0;
   27835: out<=0;
   27836: out<=1;
   27837: out<=0;
   27838: out<=0;
   27839: out<=1;
   27840: out<=1;
   27841: out<=0;
   27842: out<=0;
   27843: out<=1;
   27844: out<=0;
   27845: out<=0;
   27846: out<=0;
   27847: out<=0;
   27848: out<=1;
   27849: out<=1;
   27850: out<=0;
   27851: out<=0;
   27852: out<=0;
   27853: out<=1;
   27854: out<=0;
   27855: out<=1;
   27856: out<=0;
   27857: out<=0;
   27858: out<=0;
   27859: out<=0;
   27860: out<=0;
   27861: out<=1;
   27862: out<=1;
   27863: out<=0;
   27864: out<=1;
   27865: out<=0;
   27866: out<=1;
   27867: out<=0;
   27868: out<=1;
   27869: out<=1;
   27870: out<=0;
   27871: out<=0;
   27872: out<=0;
   27873: out<=0;
   27874: out<=1;
   27875: out<=1;
   27876: out<=0;
   27877: out<=1;
   27878: out<=0;
   27879: out<=1;
   27880: out<=0;
   27881: out<=1;
   27882: out<=1;
   27883: out<=0;
   27884: out<=0;
   27885: out<=0;
   27886: out<=0;
   27887: out<=0;
   27888: out<=1;
   27889: out<=0;
   27890: out<=1;
   27891: out<=0;
   27892: out<=0;
   27893: out<=0;
   27894: out<=1;
   27895: out<=1;
   27896: out<=0;
   27897: out<=0;
   27898: out<=0;
   27899: out<=0;
   27900: out<=1;
   27901: out<=0;
   27902: out<=0;
   27903: out<=1;
   27904: out<=1;
   27905: out<=1;
   27906: out<=1;
   27907: out<=1;
   27908: out<=1;
   27909: out<=0;
   27910: out<=0;
   27911: out<=1;
   27912: out<=0;
   27913: out<=1;
   27914: out<=0;
   27915: out<=1;
   27916: out<=0;
   27917: out<=0;
   27918: out<=1;
   27919: out<=1;
   27920: out<=1;
   27921: out<=0;
   27922: out<=0;
   27923: out<=1;
   27924: out<=0;
   27925: out<=0;
   27926: out<=0;
   27927: out<=0;
   27928: out<=1;
   27929: out<=1;
   27930: out<=0;
   27931: out<=0;
   27932: out<=0;
   27933: out<=1;
   27934: out<=0;
   27935: out<=1;
   27936: out<=0;
   27937: out<=1;
   27938: out<=0;
   27939: out<=1;
   27940: out<=1;
   27941: out<=1;
   27942: out<=0;
   27943: out<=0;
   27944: out<=1;
   27945: out<=1;
   27946: out<=1;
   27947: out<=1;
   27948: out<=0;
   27949: out<=1;
   27950: out<=1;
   27951: out<=0;
   27952: out<=0;
   27953: out<=0;
   27954: out<=1;
   27955: out<=1;
   27956: out<=0;
   27957: out<=1;
   27958: out<=0;
   27959: out<=1;
   27960: out<=0;
   27961: out<=1;
   27962: out<=1;
   27963: out<=0;
   27964: out<=0;
   27965: out<=0;
   27966: out<=0;
   27967: out<=0;
   27968: out<=0;
   27969: out<=0;
   27970: out<=0;
   27971: out<=0;
   27972: out<=0;
   27973: out<=1;
   27974: out<=1;
   27975: out<=0;
   27976: out<=1;
   27977: out<=0;
   27978: out<=1;
   27979: out<=0;
   27980: out<=1;
   27981: out<=1;
   27982: out<=0;
   27983: out<=0;
   27984: out<=1;
   27985: out<=0;
   27986: out<=0;
   27987: out<=1;
   27988: out<=0;
   27989: out<=0;
   27990: out<=0;
   27991: out<=0;
   27992: out<=1;
   27993: out<=1;
   27994: out<=0;
   27995: out<=0;
   27996: out<=0;
   27997: out<=1;
   27998: out<=0;
   27999: out<=1;
   28000: out<=0;
   28001: out<=1;
   28002: out<=0;
   28003: out<=1;
   28004: out<=1;
   28005: out<=1;
   28006: out<=0;
   28007: out<=0;
   28008: out<=1;
   28009: out<=1;
   28010: out<=1;
   28011: out<=1;
   28012: out<=0;
   28013: out<=1;
   28014: out<=1;
   28015: out<=0;
   28016: out<=1;
   28017: out<=1;
   28018: out<=0;
   28019: out<=0;
   28020: out<=1;
   28021: out<=0;
   28022: out<=1;
   28023: out<=0;
   28024: out<=1;
   28025: out<=0;
   28026: out<=0;
   28027: out<=1;
   28028: out<=1;
   28029: out<=1;
   28030: out<=1;
   28031: out<=1;
   28032: out<=0;
   28033: out<=0;
   28034: out<=0;
   28035: out<=0;
   28036: out<=0;
   28037: out<=1;
   28038: out<=1;
   28039: out<=0;
   28040: out<=1;
   28041: out<=0;
   28042: out<=1;
   28043: out<=0;
   28044: out<=1;
   28045: out<=1;
   28046: out<=0;
   28047: out<=0;
   28048: out<=1;
   28049: out<=0;
   28050: out<=0;
   28051: out<=1;
   28052: out<=0;
   28053: out<=0;
   28054: out<=0;
   28055: out<=0;
   28056: out<=1;
   28057: out<=1;
   28058: out<=0;
   28059: out<=0;
   28060: out<=0;
   28061: out<=1;
   28062: out<=0;
   28063: out<=1;
   28064: out<=1;
   28065: out<=0;
   28066: out<=1;
   28067: out<=0;
   28068: out<=0;
   28069: out<=0;
   28070: out<=1;
   28071: out<=1;
   28072: out<=0;
   28073: out<=0;
   28074: out<=0;
   28075: out<=0;
   28076: out<=1;
   28077: out<=0;
   28078: out<=0;
   28079: out<=1;
   28080: out<=0;
   28081: out<=0;
   28082: out<=1;
   28083: out<=1;
   28084: out<=0;
   28085: out<=1;
   28086: out<=0;
   28087: out<=1;
   28088: out<=0;
   28089: out<=1;
   28090: out<=1;
   28091: out<=0;
   28092: out<=0;
   28093: out<=0;
   28094: out<=0;
   28095: out<=0;
   28096: out<=1;
   28097: out<=1;
   28098: out<=1;
   28099: out<=1;
   28100: out<=1;
   28101: out<=0;
   28102: out<=0;
   28103: out<=1;
   28104: out<=0;
   28105: out<=1;
   28106: out<=0;
   28107: out<=1;
   28108: out<=0;
   28109: out<=0;
   28110: out<=1;
   28111: out<=1;
   28112: out<=1;
   28113: out<=0;
   28114: out<=0;
   28115: out<=1;
   28116: out<=0;
   28117: out<=0;
   28118: out<=0;
   28119: out<=0;
   28120: out<=1;
   28121: out<=1;
   28122: out<=0;
   28123: out<=0;
   28124: out<=0;
   28125: out<=1;
   28126: out<=0;
   28127: out<=1;
   28128: out<=1;
   28129: out<=0;
   28130: out<=1;
   28131: out<=0;
   28132: out<=0;
   28133: out<=0;
   28134: out<=1;
   28135: out<=1;
   28136: out<=0;
   28137: out<=0;
   28138: out<=0;
   28139: out<=0;
   28140: out<=1;
   28141: out<=0;
   28142: out<=0;
   28143: out<=1;
   28144: out<=1;
   28145: out<=1;
   28146: out<=0;
   28147: out<=0;
   28148: out<=1;
   28149: out<=0;
   28150: out<=1;
   28151: out<=0;
   28152: out<=1;
   28153: out<=0;
   28154: out<=0;
   28155: out<=1;
   28156: out<=1;
   28157: out<=1;
   28158: out<=1;
   28159: out<=1;
   28160: out<=1;
   28161: out<=1;
   28162: out<=0;
   28163: out<=0;
   28164: out<=1;
   28165: out<=0;
   28166: out<=1;
   28167: out<=0;
   28168: out<=1;
   28169: out<=0;
   28170: out<=0;
   28171: out<=1;
   28172: out<=1;
   28173: out<=1;
   28174: out<=1;
   28175: out<=1;
   28176: out<=1;
   28177: out<=0;
   28178: out<=1;
   28179: out<=0;
   28180: out<=0;
   28181: out<=0;
   28182: out<=1;
   28183: out<=1;
   28184: out<=0;
   28185: out<=0;
   28186: out<=0;
   28187: out<=0;
   28188: out<=1;
   28189: out<=0;
   28190: out<=0;
   28191: out<=1;
   28192: out<=1;
   28193: out<=0;
   28194: out<=0;
   28195: out<=1;
   28196: out<=0;
   28197: out<=0;
   28198: out<=0;
   28199: out<=0;
   28200: out<=1;
   28201: out<=1;
   28202: out<=0;
   28203: out<=0;
   28204: out<=0;
   28205: out<=1;
   28206: out<=0;
   28207: out<=1;
   28208: out<=1;
   28209: out<=1;
   28210: out<=1;
   28211: out<=1;
   28212: out<=1;
   28213: out<=0;
   28214: out<=0;
   28215: out<=1;
   28216: out<=0;
   28217: out<=1;
   28218: out<=0;
   28219: out<=1;
   28220: out<=0;
   28221: out<=0;
   28222: out<=1;
   28223: out<=1;
   28224: out<=0;
   28225: out<=0;
   28226: out<=1;
   28227: out<=1;
   28228: out<=0;
   28229: out<=1;
   28230: out<=0;
   28231: out<=1;
   28232: out<=0;
   28233: out<=1;
   28234: out<=1;
   28235: out<=0;
   28236: out<=0;
   28237: out<=0;
   28238: out<=0;
   28239: out<=0;
   28240: out<=1;
   28241: out<=0;
   28242: out<=1;
   28243: out<=0;
   28244: out<=0;
   28245: out<=0;
   28246: out<=1;
   28247: out<=1;
   28248: out<=0;
   28249: out<=0;
   28250: out<=0;
   28251: out<=0;
   28252: out<=1;
   28253: out<=0;
   28254: out<=0;
   28255: out<=1;
   28256: out<=1;
   28257: out<=0;
   28258: out<=0;
   28259: out<=1;
   28260: out<=0;
   28261: out<=0;
   28262: out<=0;
   28263: out<=0;
   28264: out<=1;
   28265: out<=1;
   28266: out<=0;
   28267: out<=0;
   28268: out<=0;
   28269: out<=1;
   28270: out<=0;
   28271: out<=1;
   28272: out<=0;
   28273: out<=0;
   28274: out<=0;
   28275: out<=0;
   28276: out<=0;
   28277: out<=1;
   28278: out<=1;
   28279: out<=0;
   28280: out<=1;
   28281: out<=0;
   28282: out<=1;
   28283: out<=0;
   28284: out<=1;
   28285: out<=1;
   28286: out<=0;
   28287: out<=0;
   28288: out<=1;
   28289: out<=1;
   28290: out<=0;
   28291: out<=0;
   28292: out<=1;
   28293: out<=0;
   28294: out<=1;
   28295: out<=0;
   28296: out<=1;
   28297: out<=0;
   28298: out<=0;
   28299: out<=1;
   28300: out<=1;
   28301: out<=1;
   28302: out<=1;
   28303: out<=1;
   28304: out<=0;
   28305: out<=1;
   28306: out<=0;
   28307: out<=1;
   28308: out<=1;
   28309: out<=1;
   28310: out<=0;
   28311: out<=0;
   28312: out<=1;
   28313: out<=1;
   28314: out<=1;
   28315: out<=1;
   28316: out<=0;
   28317: out<=1;
   28318: out<=1;
   28319: out<=0;
   28320: out<=1;
   28321: out<=0;
   28322: out<=0;
   28323: out<=1;
   28324: out<=0;
   28325: out<=0;
   28326: out<=0;
   28327: out<=0;
   28328: out<=1;
   28329: out<=1;
   28330: out<=0;
   28331: out<=0;
   28332: out<=0;
   28333: out<=1;
   28334: out<=0;
   28335: out<=1;
   28336: out<=0;
   28337: out<=0;
   28338: out<=0;
   28339: out<=0;
   28340: out<=0;
   28341: out<=1;
   28342: out<=1;
   28343: out<=0;
   28344: out<=1;
   28345: out<=0;
   28346: out<=1;
   28347: out<=0;
   28348: out<=1;
   28349: out<=1;
   28350: out<=0;
   28351: out<=0;
   28352: out<=0;
   28353: out<=0;
   28354: out<=1;
   28355: out<=1;
   28356: out<=0;
   28357: out<=1;
   28358: out<=0;
   28359: out<=1;
   28360: out<=0;
   28361: out<=1;
   28362: out<=1;
   28363: out<=0;
   28364: out<=0;
   28365: out<=0;
   28366: out<=0;
   28367: out<=0;
   28368: out<=0;
   28369: out<=1;
   28370: out<=0;
   28371: out<=1;
   28372: out<=1;
   28373: out<=1;
   28374: out<=0;
   28375: out<=0;
   28376: out<=1;
   28377: out<=1;
   28378: out<=1;
   28379: out<=1;
   28380: out<=0;
   28381: out<=1;
   28382: out<=1;
   28383: out<=0;
   28384: out<=1;
   28385: out<=0;
   28386: out<=0;
   28387: out<=1;
   28388: out<=0;
   28389: out<=0;
   28390: out<=0;
   28391: out<=0;
   28392: out<=1;
   28393: out<=1;
   28394: out<=0;
   28395: out<=0;
   28396: out<=0;
   28397: out<=1;
   28398: out<=0;
   28399: out<=1;
   28400: out<=1;
   28401: out<=1;
   28402: out<=1;
   28403: out<=1;
   28404: out<=1;
   28405: out<=0;
   28406: out<=0;
   28407: out<=1;
   28408: out<=0;
   28409: out<=1;
   28410: out<=0;
   28411: out<=1;
   28412: out<=0;
   28413: out<=0;
   28414: out<=1;
   28415: out<=1;
   28416: out<=1;
   28417: out<=0;
   28418: out<=1;
   28419: out<=0;
   28420: out<=0;
   28421: out<=0;
   28422: out<=1;
   28423: out<=1;
   28424: out<=0;
   28425: out<=0;
   28426: out<=0;
   28427: out<=0;
   28428: out<=1;
   28429: out<=0;
   28430: out<=0;
   28431: out<=1;
   28432: out<=0;
   28433: out<=0;
   28434: out<=1;
   28435: out<=1;
   28436: out<=0;
   28437: out<=1;
   28438: out<=0;
   28439: out<=1;
   28440: out<=0;
   28441: out<=1;
   28442: out<=1;
   28443: out<=0;
   28444: out<=0;
   28445: out<=0;
   28446: out<=0;
   28447: out<=0;
   28448: out<=0;
   28449: out<=0;
   28450: out<=0;
   28451: out<=0;
   28452: out<=0;
   28453: out<=1;
   28454: out<=1;
   28455: out<=0;
   28456: out<=1;
   28457: out<=0;
   28458: out<=1;
   28459: out<=0;
   28460: out<=1;
   28461: out<=1;
   28462: out<=0;
   28463: out<=0;
   28464: out<=1;
   28465: out<=0;
   28466: out<=0;
   28467: out<=1;
   28468: out<=0;
   28469: out<=0;
   28470: out<=0;
   28471: out<=0;
   28472: out<=1;
   28473: out<=1;
   28474: out<=0;
   28475: out<=0;
   28476: out<=0;
   28477: out<=1;
   28478: out<=0;
   28479: out<=1;
   28480: out<=1;
   28481: out<=0;
   28482: out<=1;
   28483: out<=0;
   28484: out<=0;
   28485: out<=0;
   28486: out<=1;
   28487: out<=1;
   28488: out<=0;
   28489: out<=0;
   28490: out<=0;
   28491: out<=0;
   28492: out<=1;
   28493: out<=0;
   28494: out<=0;
   28495: out<=1;
   28496: out<=1;
   28497: out<=1;
   28498: out<=0;
   28499: out<=0;
   28500: out<=1;
   28501: out<=0;
   28502: out<=1;
   28503: out<=0;
   28504: out<=1;
   28505: out<=0;
   28506: out<=0;
   28507: out<=1;
   28508: out<=1;
   28509: out<=1;
   28510: out<=1;
   28511: out<=1;
   28512: out<=1;
   28513: out<=1;
   28514: out<=1;
   28515: out<=1;
   28516: out<=1;
   28517: out<=0;
   28518: out<=0;
   28519: out<=1;
   28520: out<=0;
   28521: out<=1;
   28522: out<=0;
   28523: out<=1;
   28524: out<=0;
   28525: out<=0;
   28526: out<=1;
   28527: out<=1;
   28528: out<=1;
   28529: out<=0;
   28530: out<=0;
   28531: out<=1;
   28532: out<=0;
   28533: out<=0;
   28534: out<=0;
   28535: out<=0;
   28536: out<=1;
   28537: out<=1;
   28538: out<=0;
   28539: out<=0;
   28540: out<=0;
   28541: out<=1;
   28542: out<=0;
   28543: out<=1;
   28544: out<=0;
   28545: out<=1;
   28546: out<=0;
   28547: out<=1;
   28548: out<=1;
   28549: out<=1;
   28550: out<=0;
   28551: out<=0;
   28552: out<=1;
   28553: out<=1;
   28554: out<=1;
   28555: out<=1;
   28556: out<=0;
   28557: out<=1;
   28558: out<=1;
   28559: out<=0;
   28560: out<=0;
   28561: out<=0;
   28562: out<=1;
   28563: out<=1;
   28564: out<=0;
   28565: out<=1;
   28566: out<=0;
   28567: out<=1;
   28568: out<=0;
   28569: out<=1;
   28570: out<=1;
   28571: out<=0;
   28572: out<=0;
   28573: out<=0;
   28574: out<=0;
   28575: out<=0;
   28576: out<=1;
   28577: out<=1;
   28578: out<=1;
   28579: out<=1;
   28580: out<=1;
   28581: out<=0;
   28582: out<=0;
   28583: out<=1;
   28584: out<=0;
   28585: out<=1;
   28586: out<=0;
   28587: out<=1;
   28588: out<=0;
   28589: out<=0;
   28590: out<=1;
   28591: out<=1;
   28592: out<=1;
   28593: out<=0;
   28594: out<=0;
   28595: out<=1;
   28596: out<=0;
   28597: out<=0;
   28598: out<=0;
   28599: out<=0;
   28600: out<=1;
   28601: out<=1;
   28602: out<=0;
   28603: out<=0;
   28604: out<=0;
   28605: out<=1;
   28606: out<=0;
   28607: out<=1;
   28608: out<=0;
   28609: out<=1;
   28610: out<=0;
   28611: out<=1;
   28612: out<=1;
   28613: out<=1;
   28614: out<=0;
   28615: out<=0;
   28616: out<=1;
   28617: out<=1;
   28618: out<=1;
   28619: out<=1;
   28620: out<=0;
   28621: out<=1;
   28622: out<=1;
   28623: out<=0;
   28624: out<=1;
   28625: out<=1;
   28626: out<=0;
   28627: out<=0;
   28628: out<=1;
   28629: out<=0;
   28630: out<=1;
   28631: out<=0;
   28632: out<=1;
   28633: out<=0;
   28634: out<=0;
   28635: out<=1;
   28636: out<=1;
   28637: out<=1;
   28638: out<=1;
   28639: out<=1;
   28640: out<=0;
   28641: out<=0;
   28642: out<=0;
   28643: out<=0;
   28644: out<=0;
   28645: out<=1;
   28646: out<=1;
   28647: out<=0;
   28648: out<=1;
   28649: out<=0;
   28650: out<=1;
   28651: out<=0;
   28652: out<=1;
   28653: out<=1;
   28654: out<=0;
   28655: out<=0;
   28656: out<=1;
   28657: out<=0;
   28658: out<=0;
   28659: out<=1;
   28660: out<=0;
   28661: out<=0;
   28662: out<=0;
   28663: out<=0;
   28664: out<=1;
   28665: out<=1;
   28666: out<=0;
   28667: out<=0;
   28668: out<=0;
   28669: out<=1;
   28670: out<=0;
   28671: out<=1;
   28672: out<=0;
   28673: out<=1;
   28674: out<=0;
   28675: out<=1;
   28676: out<=0;
   28677: out<=0;
   28678: out<=1;
   28679: out<=1;
   28680: out<=1;
   28681: out<=1;
   28682: out<=1;
   28683: out<=1;
   28684: out<=1;
   28685: out<=0;
   28686: out<=0;
   28687: out<=1;
   28688: out<=1;
   28689: out<=1;
   28690: out<=0;
   28691: out<=0;
   28692: out<=0;
   28693: out<=1;
   28694: out<=0;
   28695: out<=1;
   28696: out<=1;
   28697: out<=0;
   28698: out<=0;
   28699: out<=1;
   28700: out<=0;
   28701: out<=0;
   28702: out<=0;
   28703: out<=0;
   28704: out<=0;
   28705: out<=0;
   28706: out<=0;
   28707: out<=0;
   28708: out<=1;
   28709: out<=0;
   28710: out<=0;
   28711: out<=1;
   28712: out<=1;
   28713: out<=0;
   28714: out<=1;
   28715: out<=0;
   28716: out<=0;
   28717: out<=0;
   28718: out<=1;
   28719: out<=1;
   28720: out<=1;
   28721: out<=0;
   28722: out<=0;
   28723: out<=1;
   28724: out<=1;
   28725: out<=1;
   28726: out<=1;
   28727: out<=1;
   28728: out<=1;
   28729: out<=1;
   28730: out<=0;
   28731: out<=0;
   28732: out<=1;
   28733: out<=0;
   28734: out<=1;
   28735: out<=0;
   28736: out<=0;
   28737: out<=1;
   28738: out<=0;
   28739: out<=1;
   28740: out<=0;
   28741: out<=0;
   28742: out<=1;
   28743: out<=1;
   28744: out<=1;
   28745: out<=1;
   28746: out<=1;
   28747: out<=1;
   28748: out<=1;
   28749: out<=0;
   28750: out<=0;
   28751: out<=1;
   28752: out<=0;
   28753: out<=0;
   28754: out<=1;
   28755: out<=1;
   28756: out<=1;
   28757: out<=0;
   28758: out<=1;
   28759: out<=0;
   28760: out<=0;
   28761: out<=1;
   28762: out<=1;
   28763: out<=0;
   28764: out<=1;
   28765: out<=1;
   28766: out<=1;
   28767: out<=1;
   28768: out<=1;
   28769: out<=1;
   28770: out<=1;
   28771: out<=1;
   28772: out<=0;
   28773: out<=1;
   28774: out<=1;
   28775: out<=0;
   28776: out<=0;
   28777: out<=1;
   28778: out<=0;
   28779: out<=1;
   28780: out<=1;
   28781: out<=1;
   28782: out<=0;
   28783: out<=0;
   28784: out<=1;
   28785: out<=0;
   28786: out<=0;
   28787: out<=1;
   28788: out<=1;
   28789: out<=1;
   28790: out<=1;
   28791: out<=1;
   28792: out<=1;
   28793: out<=1;
   28794: out<=0;
   28795: out<=0;
   28796: out<=1;
   28797: out<=0;
   28798: out<=1;
   28799: out<=0;
   28800: out<=1;
   28801: out<=0;
   28802: out<=1;
   28803: out<=0;
   28804: out<=1;
   28805: out<=1;
   28806: out<=0;
   28807: out<=0;
   28808: out<=0;
   28809: out<=0;
   28810: out<=0;
   28811: out<=0;
   28812: out<=0;
   28813: out<=1;
   28814: out<=1;
   28815: out<=0;
   28816: out<=1;
   28817: out<=1;
   28818: out<=0;
   28819: out<=0;
   28820: out<=0;
   28821: out<=1;
   28822: out<=0;
   28823: out<=1;
   28824: out<=1;
   28825: out<=0;
   28826: out<=0;
   28827: out<=1;
   28828: out<=0;
   28829: out<=0;
   28830: out<=0;
   28831: out<=0;
   28832: out<=1;
   28833: out<=1;
   28834: out<=1;
   28835: out<=1;
   28836: out<=0;
   28837: out<=1;
   28838: out<=1;
   28839: out<=0;
   28840: out<=0;
   28841: out<=1;
   28842: out<=0;
   28843: out<=1;
   28844: out<=1;
   28845: out<=1;
   28846: out<=0;
   28847: out<=0;
   28848: out<=1;
   28849: out<=0;
   28850: out<=0;
   28851: out<=1;
   28852: out<=1;
   28853: out<=1;
   28854: out<=1;
   28855: out<=1;
   28856: out<=1;
   28857: out<=1;
   28858: out<=0;
   28859: out<=0;
   28860: out<=1;
   28861: out<=0;
   28862: out<=1;
   28863: out<=0;
   28864: out<=1;
   28865: out<=0;
   28866: out<=1;
   28867: out<=0;
   28868: out<=1;
   28869: out<=1;
   28870: out<=0;
   28871: out<=0;
   28872: out<=0;
   28873: out<=0;
   28874: out<=0;
   28875: out<=0;
   28876: out<=0;
   28877: out<=1;
   28878: out<=1;
   28879: out<=0;
   28880: out<=0;
   28881: out<=0;
   28882: out<=1;
   28883: out<=1;
   28884: out<=1;
   28885: out<=0;
   28886: out<=1;
   28887: out<=0;
   28888: out<=0;
   28889: out<=1;
   28890: out<=1;
   28891: out<=0;
   28892: out<=1;
   28893: out<=1;
   28894: out<=1;
   28895: out<=1;
   28896: out<=0;
   28897: out<=0;
   28898: out<=0;
   28899: out<=0;
   28900: out<=1;
   28901: out<=0;
   28902: out<=0;
   28903: out<=1;
   28904: out<=1;
   28905: out<=0;
   28906: out<=1;
   28907: out<=0;
   28908: out<=0;
   28909: out<=0;
   28910: out<=1;
   28911: out<=1;
   28912: out<=1;
   28913: out<=0;
   28914: out<=0;
   28915: out<=1;
   28916: out<=1;
   28917: out<=1;
   28918: out<=1;
   28919: out<=1;
   28920: out<=1;
   28921: out<=1;
   28922: out<=0;
   28923: out<=0;
   28924: out<=1;
   28925: out<=0;
   28926: out<=1;
   28927: out<=0;
   28928: out<=0;
   28929: out<=0;
   28930: out<=1;
   28931: out<=1;
   28932: out<=1;
   28933: out<=0;
   28934: out<=1;
   28935: out<=0;
   28936: out<=0;
   28937: out<=1;
   28938: out<=1;
   28939: out<=0;
   28940: out<=1;
   28941: out<=1;
   28942: out<=1;
   28943: out<=1;
   28944: out<=0;
   28945: out<=1;
   28946: out<=0;
   28947: out<=1;
   28948: out<=0;
   28949: out<=0;
   28950: out<=1;
   28951: out<=1;
   28952: out<=1;
   28953: out<=1;
   28954: out<=1;
   28955: out<=1;
   28956: out<=1;
   28957: out<=0;
   28958: out<=0;
   28959: out<=1;
   28960: out<=1;
   28961: out<=0;
   28962: out<=0;
   28963: out<=1;
   28964: out<=1;
   28965: out<=1;
   28966: out<=1;
   28967: out<=1;
   28968: out<=1;
   28969: out<=1;
   28970: out<=0;
   28971: out<=0;
   28972: out<=1;
   28973: out<=0;
   28974: out<=1;
   28975: out<=0;
   28976: out<=1;
   28977: out<=1;
   28978: out<=1;
   28979: out<=1;
   28980: out<=0;
   28981: out<=1;
   28982: out<=1;
   28983: out<=0;
   28984: out<=0;
   28985: out<=1;
   28986: out<=0;
   28987: out<=1;
   28988: out<=1;
   28989: out<=1;
   28990: out<=0;
   28991: out<=0;
   28992: out<=1;
   28993: out<=1;
   28994: out<=0;
   28995: out<=0;
   28996: out<=0;
   28997: out<=1;
   28998: out<=0;
   28999: out<=1;
   29000: out<=1;
   29001: out<=0;
   29002: out<=0;
   29003: out<=1;
   29004: out<=0;
   29005: out<=0;
   29006: out<=0;
   29007: out<=0;
   29008: out<=0;
   29009: out<=1;
   29010: out<=0;
   29011: out<=1;
   29012: out<=0;
   29013: out<=0;
   29014: out<=1;
   29015: out<=1;
   29016: out<=1;
   29017: out<=1;
   29018: out<=1;
   29019: out<=1;
   29020: out<=1;
   29021: out<=0;
   29022: out<=0;
   29023: out<=1;
   29024: out<=1;
   29025: out<=0;
   29026: out<=0;
   29027: out<=1;
   29028: out<=1;
   29029: out<=1;
   29030: out<=1;
   29031: out<=1;
   29032: out<=1;
   29033: out<=1;
   29034: out<=0;
   29035: out<=0;
   29036: out<=1;
   29037: out<=0;
   29038: out<=1;
   29039: out<=0;
   29040: out<=0;
   29041: out<=0;
   29042: out<=0;
   29043: out<=0;
   29044: out<=1;
   29045: out<=0;
   29046: out<=0;
   29047: out<=1;
   29048: out<=1;
   29049: out<=0;
   29050: out<=1;
   29051: out<=0;
   29052: out<=0;
   29053: out<=0;
   29054: out<=1;
   29055: out<=1;
   29056: out<=0;
   29057: out<=0;
   29058: out<=1;
   29059: out<=1;
   29060: out<=1;
   29061: out<=0;
   29062: out<=1;
   29063: out<=0;
   29064: out<=0;
   29065: out<=1;
   29066: out<=1;
   29067: out<=0;
   29068: out<=1;
   29069: out<=1;
   29070: out<=1;
   29071: out<=1;
   29072: out<=1;
   29073: out<=0;
   29074: out<=1;
   29075: out<=0;
   29076: out<=1;
   29077: out<=1;
   29078: out<=0;
   29079: out<=0;
   29080: out<=0;
   29081: out<=0;
   29082: out<=0;
   29083: out<=0;
   29084: out<=0;
   29085: out<=1;
   29086: out<=1;
   29087: out<=0;
   29088: out<=1;
   29089: out<=0;
   29090: out<=0;
   29091: out<=1;
   29092: out<=1;
   29093: out<=1;
   29094: out<=1;
   29095: out<=1;
   29096: out<=1;
   29097: out<=1;
   29098: out<=0;
   29099: out<=0;
   29100: out<=1;
   29101: out<=0;
   29102: out<=1;
   29103: out<=0;
   29104: out<=0;
   29105: out<=0;
   29106: out<=0;
   29107: out<=0;
   29108: out<=1;
   29109: out<=0;
   29110: out<=0;
   29111: out<=1;
   29112: out<=1;
   29113: out<=0;
   29114: out<=1;
   29115: out<=0;
   29116: out<=0;
   29117: out<=0;
   29118: out<=1;
   29119: out<=1;
   29120: out<=1;
   29121: out<=1;
   29122: out<=0;
   29123: out<=0;
   29124: out<=0;
   29125: out<=1;
   29126: out<=0;
   29127: out<=1;
   29128: out<=1;
   29129: out<=0;
   29130: out<=0;
   29131: out<=1;
   29132: out<=0;
   29133: out<=0;
   29134: out<=0;
   29135: out<=0;
   29136: out<=1;
   29137: out<=0;
   29138: out<=1;
   29139: out<=0;
   29140: out<=1;
   29141: out<=1;
   29142: out<=0;
   29143: out<=0;
   29144: out<=0;
   29145: out<=0;
   29146: out<=0;
   29147: out<=0;
   29148: out<=0;
   29149: out<=1;
   29150: out<=1;
   29151: out<=0;
   29152: out<=1;
   29153: out<=0;
   29154: out<=0;
   29155: out<=1;
   29156: out<=1;
   29157: out<=1;
   29158: out<=1;
   29159: out<=1;
   29160: out<=1;
   29161: out<=1;
   29162: out<=0;
   29163: out<=0;
   29164: out<=1;
   29165: out<=0;
   29166: out<=1;
   29167: out<=0;
   29168: out<=1;
   29169: out<=1;
   29170: out<=1;
   29171: out<=1;
   29172: out<=0;
   29173: out<=1;
   29174: out<=1;
   29175: out<=0;
   29176: out<=0;
   29177: out<=1;
   29178: out<=0;
   29179: out<=1;
   29180: out<=1;
   29181: out<=1;
   29182: out<=0;
   29183: out<=0;
   29184: out<=1;
   29185: out<=1;
   29186: out<=1;
   29187: out<=1;
   29188: out<=0;
   29189: out<=1;
   29190: out<=1;
   29191: out<=0;
   29192: out<=0;
   29193: out<=1;
   29194: out<=0;
   29195: out<=1;
   29196: out<=1;
   29197: out<=1;
   29198: out<=0;
   29199: out<=0;
   29200: out<=1;
   29201: out<=0;
   29202: out<=0;
   29203: out<=1;
   29204: out<=1;
   29205: out<=1;
   29206: out<=1;
   29207: out<=1;
   29208: out<=1;
   29209: out<=1;
   29210: out<=0;
   29211: out<=0;
   29212: out<=1;
   29213: out<=0;
   29214: out<=1;
   29215: out<=0;
   29216: out<=1;
   29217: out<=0;
   29218: out<=1;
   29219: out<=0;
   29220: out<=1;
   29221: out<=1;
   29222: out<=0;
   29223: out<=0;
   29224: out<=0;
   29225: out<=0;
   29226: out<=0;
   29227: out<=0;
   29228: out<=0;
   29229: out<=1;
   29230: out<=1;
   29231: out<=0;
   29232: out<=1;
   29233: out<=1;
   29234: out<=0;
   29235: out<=0;
   29236: out<=0;
   29237: out<=1;
   29238: out<=0;
   29239: out<=1;
   29240: out<=1;
   29241: out<=0;
   29242: out<=0;
   29243: out<=1;
   29244: out<=0;
   29245: out<=0;
   29246: out<=0;
   29247: out<=0;
   29248: out<=0;
   29249: out<=0;
   29250: out<=0;
   29251: out<=0;
   29252: out<=1;
   29253: out<=0;
   29254: out<=0;
   29255: out<=1;
   29256: out<=1;
   29257: out<=0;
   29258: out<=1;
   29259: out<=0;
   29260: out<=0;
   29261: out<=0;
   29262: out<=1;
   29263: out<=1;
   29264: out<=1;
   29265: out<=0;
   29266: out<=0;
   29267: out<=1;
   29268: out<=1;
   29269: out<=1;
   29270: out<=1;
   29271: out<=1;
   29272: out<=1;
   29273: out<=1;
   29274: out<=0;
   29275: out<=0;
   29276: out<=1;
   29277: out<=0;
   29278: out<=1;
   29279: out<=0;
   29280: out<=1;
   29281: out<=0;
   29282: out<=1;
   29283: out<=0;
   29284: out<=1;
   29285: out<=1;
   29286: out<=0;
   29287: out<=0;
   29288: out<=0;
   29289: out<=0;
   29290: out<=0;
   29291: out<=0;
   29292: out<=0;
   29293: out<=1;
   29294: out<=1;
   29295: out<=0;
   29296: out<=0;
   29297: out<=0;
   29298: out<=1;
   29299: out<=1;
   29300: out<=1;
   29301: out<=0;
   29302: out<=1;
   29303: out<=0;
   29304: out<=0;
   29305: out<=1;
   29306: out<=1;
   29307: out<=0;
   29308: out<=1;
   29309: out<=1;
   29310: out<=1;
   29311: out<=1;
   29312: out<=0;
   29313: out<=0;
   29314: out<=0;
   29315: out<=0;
   29316: out<=1;
   29317: out<=0;
   29318: out<=0;
   29319: out<=1;
   29320: out<=1;
   29321: out<=0;
   29322: out<=1;
   29323: out<=0;
   29324: out<=0;
   29325: out<=0;
   29326: out<=1;
   29327: out<=1;
   29328: out<=1;
   29329: out<=0;
   29330: out<=0;
   29331: out<=1;
   29332: out<=1;
   29333: out<=1;
   29334: out<=1;
   29335: out<=1;
   29336: out<=1;
   29337: out<=1;
   29338: out<=0;
   29339: out<=0;
   29340: out<=1;
   29341: out<=0;
   29342: out<=1;
   29343: out<=0;
   29344: out<=0;
   29345: out<=1;
   29346: out<=0;
   29347: out<=1;
   29348: out<=0;
   29349: out<=0;
   29350: out<=1;
   29351: out<=1;
   29352: out<=1;
   29353: out<=1;
   29354: out<=1;
   29355: out<=1;
   29356: out<=1;
   29357: out<=0;
   29358: out<=0;
   29359: out<=1;
   29360: out<=1;
   29361: out<=1;
   29362: out<=0;
   29363: out<=0;
   29364: out<=0;
   29365: out<=1;
   29366: out<=0;
   29367: out<=1;
   29368: out<=1;
   29369: out<=0;
   29370: out<=0;
   29371: out<=1;
   29372: out<=0;
   29373: out<=0;
   29374: out<=0;
   29375: out<=0;
   29376: out<=1;
   29377: out<=1;
   29378: out<=1;
   29379: out<=1;
   29380: out<=0;
   29381: out<=1;
   29382: out<=1;
   29383: out<=0;
   29384: out<=0;
   29385: out<=1;
   29386: out<=0;
   29387: out<=1;
   29388: out<=1;
   29389: out<=1;
   29390: out<=0;
   29391: out<=0;
   29392: out<=1;
   29393: out<=0;
   29394: out<=0;
   29395: out<=1;
   29396: out<=1;
   29397: out<=1;
   29398: out<=1;
   29399: out<=1;
   29400: out<=1;
   29401: out<=1;
   29402: out<=0;
   29403: out<=0;
   29404: out<=1;
   29405: out<=0;
   29406: out<=1;
   29407: out<=0;
   29408: out<=0;
   29409: out<=1;
   29410: out<=0;
   29411: out<=1;
   29412: out<=0;
   29413: out<=0;
   29414: out<=1;
   29415: out<=1;
   29416: out<=1;
   29417: out<=1;
   29418: out<=1;
   29419: out<=1;
   29420: out<=1;
   29421: out<=0;
   29422: out<=0;
   29423: out<=1;
   29424: out<=0;
   29425: out<=0;
   29426: out<=1;
   29427: out<=1;
   29428: out<=1;
   29429: out<=0;
   29430: out<=1;
   29431: out<=0;
   29432: out<=0;
   29433: out<=1;
   29434: out<=1;
   29435: out<=0;
   29436: out<=1;
   29437: out<=1;
   29438: out<=1;
   29439: out<=1;
   29440: out<=1;
   29441: out<=0;
   29442: out<=0;
   29443: out<=1;
   29444: out<=1;
   29445: out<=1;
   29446: out<=1;
   29447: out<=1;
   29448: out<=1;
   29449: out<=1;
   29450: out<=0;
   29451: out<=0;
   29452: out<=1;
   29453: out<=0;
   29454: out<=1;
   29455: out<=0;
   29456: out<=0;
   29457: out<=0;
   29458: out<=0;
   29459: out<=0;
   29460: out<=1;
   29461: out<=0;
   29462: out<=0;
   29463: out<=1;
   29464: out<=1;
   29465: out<=0;
   29466: out<=1;
   29467: out<=0;
   29468: out<=0;
   29469: out<=0;
   29470: out<=1;
   29471: out<=1;
   29472: out<=0;
   29473: out<=0;
   29474: out<=1;
   29475: out<=1;
   29476: out<=1;
   29477: out<=0;
   29478: out<=1;
   29479: out<=0;
   29480: out<=0;
   29481: out<=1;
   29482: out<=1;
   29483: out<=0;
   29484: out<=1;
   29485: out<=1;
   29486: out<=1;
   29487: out<=1;
   29488: out<=1;
   29489: out<=0;
   29490: out<=1;
   29491: out<=0;
   29492: out<=1;
   29493: out<=1;
   29494: out<=0;
   29495: out<=0;
   29496: out<=0;
   29497: out<=0;
   29498: out<=0;
   29499: out<=0;
   29500: out<=0;
   29501: out<=1;
   29502: out<=1;
   29503: out<=0;
   29504: out<=1;
   29505: out<=0;
   29506: out<=0;
   29507: out<=1;
   29508: out<=1;
   29509: out<=1;
   29510: out<=1;
   29511: out<=1;
   29512: out<=1;
   29513: out<=1;
   29514: out<=0;
   29515: out<=0;
   29516: out<=1;
   29517: out<=0;
   29518: out<=1;
   29519: out<=0;
   29520: out<=1;
   29521: out<=1;
   29522: out<=1;
   29523: out<=1;
   29524: out<=0;
   29525: out<=1;
   29526: out<=1;
   29527: out<=0;
   29528: out<=0;
   29529: out<=1;
   29530: out<=0;
   29531: out<=1;
   29532: out<=1;
   29533: out<=1;
   29534: out<=0;
   29535: out<=0;
   29536: out<=1;
   29537: out<=1;
   29538: out<=0;
   29539: out<=0;
   29540: out<=0;
   29541: out<=1;
   29542: out<=0;
   29543: out<=1;
   29544: out<=1;
   29545: out<=0;
   29546: out<=0;
   29547: out<=1;
   29548: out<=0;
   29549: out<=0;
   29550: out<=0;
   29551: out<=0;
   29552: out<=1;
   29553: out<=0;
   29554: out<=1;
   29555: out<=0;
   29556: out<=1;
   29557: out<=1;
   29558: out<=0;
   29559: out<=0;
   29560: out<=0;
   29561: out<=0;
   29562: out<=0;
   29563: out<=0;
   29564: out<=0;
   29565: out<=1;
   29566: out<=1;
   29567: out<=0;
   29568: out<=1;
   29569: out<=0;
   29570: out<=0;
   29571: out<=1;
   29572: out<=1;
   29573: out<=1;
   29574: out<=1;
   29575: out<=1;
   29576: out<=1;
   29577: out<=1;
   29578: out<=0;
   29579: out<=0;
   29580: out<=1;
   29581: out<=0;
   29582: out<=1;
   29583: out<=0;
   29584: out<=1;
   29585: out<=1;
   29586: out<=1;
   29587: out<=1;
   29588: out<=0;
   29589: out<=1;
   29590: out<=1;
   29591: out<=0;
   29592: out<=0;
   29593: out<=1;
   29594: out<=0;
   29595: out<=1;
   29596: out<=1;
   29597: out<=1;
   29598: out<=0;
   29599: out<=0;
   29600: out<=0;
   29601: out<=0;
   29602: out<=1;
   29603: out<=1;
   29604: out<=1;
   29605: out<=0;
   29606: out<=1;
   29607: out<=0;
   29608: out<=0;
   29609: out<=1;
   29610: out<=1;
   29611: out<=0;
   29612: out<=1;
   29613: out<=1;
   29614: out<=1;
   29615: out<=1;
   29616: out<=0;
   29617: out<=1;
   29618: out<=0;
   29619: out<=1;
   29620: out<=0;
   29621: out<=0;
   29622: out<=1;
   29623: out<=1;
   29624: out<=1;
   29625: out<=1;
   29626: out<=1;
   29627: out<=1;
   29628: out<=1;
   29629: out<=0;
   29630: out<=0;
   29631: out<=1;
   29632: out<=1;
   29633: out<=0;
   29634: out<=0;
   29635: out<=1;
   29636: out<=1;
   29637: out<=1;
   29638: out<=1;
   29639: out<=1;
   29640: out<=1;
   29641: out<=1;
   29642: out<=0;
   29643: out<=0;
   29644: out<=1;
   29645: out<=0;
   29646: out<=1;
   29647: out<=0;
   29648: out<=0;
   29649: out<=0;
   29650: out<=0;
   29651: out<=0;
   29652: out<=1;
   29653: out<=0;
   29654: out<=0;
   29655: out<=1;
   29656: out<=1;
   29657: out<=0;
   29658: out<=1;
   29659: out<=0;
   29660: out<=0;
   29661: out<=0;
   29662: out<=1;
   29663: out<=1;
   29664: out<=1;
   29665: out<=1;
   29666: out<=0;
   29667: out<=0;
   29668: out<=0;
   29669: out<=1;
   29670: out<=0;
   29671: out<=1;
   29672: out<=1;
   29673: out<=0;
   29674: out<=0;
   29675: out<=1;
   29676: out<=0;
   29677: out<=0;
   29678: out<=0;
   29679: out<=0;
   29680: out<=0;
   29681: out<=1;
   29682: out<=0;
   29683: out<=1;
   29684: out<=0;
   29685: out<=0;
   29686: out<=1;
   29687: out<=1;
   29688: out<=1;
   29689: out<=1;
   29690: out<=1;
   29691: out<=1;
   29692: out<=1;
   29693: out<=0;
   29694: out<=0;
   29695: out<=1;
   29696: out<=0;
   29697: out<=0;
   29698: out<=1;
   29699: out<=1;
   29700: out<=0;
   29701: out<=1;
   29702: out<=0;
   29703: out<=1;
   29704: out<=1;
   29705: out<=0;
   29706: out<=0;
   29707: out<=1;
   29708: out<=1;
   29709: out<=1;
   29710: out<=1;
   29711: out<=1;
   29712: out<=1;
   29713: out<=0;
   29714: out<=1;
   29715: out<=0;
   29716: out<=0;
   29717: out<=0;
   29718: out<=1;
   29719: out<=1;
   29720: out<=1;
   29721: out<=1;
   29722: out<=1;
   29723: out<=1;
   29724: out<=0;
   29725: out<=1;
   29726: out<=1;
   29727: out<=0;
   29728: out<=0;
   29729: out<=1;
   29730: out<=1;
   29731: out<=0;
   29732: out<=1;
   29733: out<=1;
   29734: out<=1;
   29735: out<=1;
   29736: out<=1;
   29737: out<=1;
   29738: out<=0;
   29739: out<=0;
   29740: out<=0;
   29741: out<=1;
   29742: out<=0;
   29743: out<=1;
   29744: out<=1;
   29745: out<=1;
   29746: out<=1;
   29747: out<=1;
   29748: out<=1;
   29749: out<=0;
   29750: out<=0;
   29751: out<=1;
   29752: out<=1;
   29753: out<=0;
   29754: out<=1;
   29755: out<=0;
   29756: out<=1;
   29757: out<=1;
   29758: out<=0;
   29759: out<=0;
   29760: out<=1;
   29761: out<=1;
   29762: out<=0;
   29763: out<=0;
   29764: out<=1;
   29765: out<=0;
   29766: out<=1;
   29767: out<=0;
   29768: out<=0;
   29769: out<=1;
   29770: out<=1;
   29771: out<=0;
   29772: out<=0;
   29773: out<=0;
   29774: out<=0;
   29775: out<=0;
   29776: out<=1;
   29777: out<=0;
   29778: out<=1;
   29779: out<=0;
   29780: out<=0;
   29781: out<=0;
   29782: out<=1;
   29783: out<=1;
   29784: out<=1;
   29785: out<=1;
   29786: out<=1;
   29787: out<=1;
   29788: out<=0;
   29789: out<=1;
   29790: out<=1;
   29791: out<=0;
   29792: out<=0;
   29793: out<=1;
   29794: out<=1;
   29795: out<=0;
   29796: out<=1;
   29797: out<=1;
   29798: out<=1;
   29799: out<=1;
   29800: out<=1;
   29801: out<=1;
   29802: out<=0;
   29803: out<=0;
   29804: out<=0;
   29805: out<=1;
   29806: out<=0;
   29807: out<=1;
   29808: out<=0;
   29809: out<=0;
   29810: out<=0;
   29811: out<=0;
   29812: out<=0;
   29813: out<=1;
   29814: out<=1;
   29815: out<=0;
   29816: out<=0;
   29817: out<=1;
   29818: out<=0;
   29819: out<=1;
   29820: out<=0;
   29821: out<=0;
   29822: out<=1;
   29823: out<=1;
   29824: out<=0;
   29825: out<=0;
   29826: out<=1;
   29827: out<=1;
   29828: out<=0;
   29829: out<=1;
   29830: out<=0;
   29831: out<=1;
   29832: out<=1;
   29833: out<=0;
   29834: out<=0;
   29835: out<=1;
   29836: out<=1;
   29837: out<=1;
   29838: out<=1;
   29839: out<=1;
   29840: out<=0;
   29841: out<=1;
   29842: out<=0;
   29843: out<=1;
   29844: out<=1;
   29845: out<=1;
   29846: out<=0;
   29847: out<=0;
   29848: out<=0;
   29849: out<=0;
   29850: out<=0;
   29851: out<=0;
   29852: out<=1;
   29853: out<=0;
   29854: out<=0;
   29855: out<=1;
   29856: out<=0;
   29857: out<=1;
   29858: out<=1;
   29859: out<=0;
   29860: out<=1;
   29861: out<=1;
   29862: out<=1;
   29863: out<=1;
   29864: out<=1;
   29865: out<=1;
   29866: out<=0;
   29867: out<=0;
   29868: out<=0;
   29869: out<=1;
   29870: out<=0;
   29871: out<=1;
   29872: out<=0;
   29873: out<=0;
   29874: out<=0;
   29875: out<=0;
   29876: out<=0;
   29877: out<=1;
   29878: out<=1;
   29879: out<=0;
   29880: out<=0;
   29881: out<=1;
   29882: out<=0;
   29883: out<=1;
   29884: out<=0;
   29885: out<=0;
   29886: out<=1;
   29887: out<=1;
   29888: out<=1;
   29889: out<=1;
   29890: out<=0;
   29891: out<=0;
   29892: out<=1;
   29893: out<=0;
   29894: out<=1;
   29895: out<=0;
   29896: out<=0;
   29897: out<=1;
   29898: out<=1;
   29899: out<=0;
   29900: out<=0;
   29901: out<=0;
   29902: out<=0;
   29903: out<=0;
   29904: out<=0;
   29905: out<=1;
   29906: out<=0;
   29907: out<=1;
   29908: out<=1;
   29909: out<=1;
   29910: out<=0;
   29911: out<=0;
   29912: out<=0;
   29913: out<=0;
   29914: out<=0;
   29915: out<=0;
   29916: out<=1;
   29917: out<=0;
   29918: out<=0;
   29919: out<=1;
   29920: out<=0;
   29921: out<=1;
   29922: out<=1;
   29923: out<=0;
   29924: out<=1;
   29925: out<=1;
   29926: out<=1;
   29927: out<=1;
   29928: out<=1;
   29929: out<=1;
   29930: out<=0;
   29931: out<=0;
   29932: out<=0;
   29933: out<=1;
   29934: out<=0;
   29935: out<=1;
   29936: out<=1;
   29937: out<=1;
   29938: out<=1;
   29939: out<=1;
   29940: out<=1;
   29941: out<=0;
   29942: out<=0;
   29943: out<=1;
   29944: out<=1;
   29945: out<=0;
   29946: out<=1;
   29947: out<=0;
   29948: out<=1;
   29949: out<=1;
   29950: out<=0;
   29951: out<=0;
   29952: out<=1;
   29953: out<=0;
   29954: out<=1;
   29955: out<=0;
   29956: out<=0;
   29957: out<=0;
   29958: out<=1;
   29959: out<=1;
   29960: out<=1;
   29961: out<=1;
   29962: out<=1;
   29963: out<=1;
   29964: out<=0;
   29965: out<=1;
   29966: out<=1;
   29967: out<=0;
   29968: out<=1;
   29969: out<=1;
   29970: out<=0;
   29971: out<=0;
   29972: out<=1;
   29973: out<=0;
   29974: out<=1;
   29975: out<=0;
   29976: out<=0;
   29977: out<=1;
   29978: out<=1;
   29979: out<=0;
   29980: out<=0;
   29981: out<=0;
   29982: out<=0;
   29983: out<=0;
   29984: out<=0;
   29985: out<=0;
   29986: out<=0;
   29987: out<=0;
   29988: out<=0;
   29989: out<=1;
   29990: out<=1;
   29991: out<=0;
   29992: out<=0;
   29993: out<=1;
   29994: out<=0;
   29995: out<=1;
   29996: out<=0;
   29997: out<=0;
   29998: out<=1;
   29999: out<=1;
   30000: out<=0;
   30001: out<=1;
   30002: out<=1;
   30003: out<=0;
   30004: out<=1;
   30005: out<=1;
   30006: out<=1;
   30007: out<=1;
   30008: out<=1;
   30009: out<=1;
   30010: out<=0;
   30011: out<=0;
   30012: out<=0;
   30013: out<=1;
   30014: out<=0;
   30015: out<=1;
   30016: out<=1;
   30017: out<=0;
   30018: out<=1;
   30019: out<=0;
   30020: out<=0;
   30021: out<=0;
   30022: out<=1;
   30023: out<=1;
   30024: out<=1;
   30025: out<=1;
   30026: out<=1;
   30027: out<=1;
   30028: out<=0;
   30029: out<=1;
   30030: out<=1;
   30031: out<=0;
   30032: out<=0;
   30033: out<=0;
   30034: out<=1;
   30035: out<=1;
   30036: out<=0;
   30037: out<=1;
   30038: out<=0;
   30039: out<=1;
   30040: out<=1;
   30041: out<=0;
   30042: out<=0;
   30043: out<=1;
   30044: out<=1;
   30045: out<=1;
   30046: out<=1;
   30047: out<=1;
   30048: out<=1;
   30049: out<=1;
   30050: out<=1;
   30051: out<=1;
   30052: out<=1;
   30053: out<=0;
   30054: out<=0;
   30055: out<=1;
   30056: out<=1;
   30057: out<=0;
   30058: out<=1;
   30059: out<=0;
   30060: out<=1;
   30061: out<=1;
   30062: out<=0;
   30063: out<=0;
   30064: out<=0;
   30065: out<=1;
   30066: out<=1;
   30067: out<=0;
   30068: out<=1;
   30069: out<=1;
   30070: out<=1;
   30071: out<=1;
   30072: out<=1;
   30073: out<=1;
   30074: out<=0;
   30075: out<=0;
   30076: out<=0;
   30077: out<=1;
   30078: out<=0;
   30079: out<=1;
   30080: out<=0;
   30081: out<=1;
   30082: out<=0;
   30083: out<=1;
   30084: out<=1;
   30085: out<=1;
   30086: out<=0;
   30087: out<=0;
   30088: out<=0;
   30089: out<=0;
   30090: out<=0;
   30091: out<=0;
   30092: out<=1;
   30093: out<=0;
   30094: out<=0;
   30095: out<=1;
   30096: out<=1;
   30097: out<=1;
   30098: out<=0;
   30099: out<=0;
   30100: out<=1;
   30101: out<=0;
   30102: out<=1;
   30103: out<=0;
   30104: out<=0;
   30105: out<=1;
   30106: out<=1;
   30107: out<=0;
   30108: out<=0;
   30109: out<=0;
   30110: out<=0;
   30111: out<=0;
   30112: out<=1;
   30113: out<=1;
   30114: out<=1;
   30115: out<=1;
   30116: out<=1;
   30117: out<=0;
   30118: out<=0;
   30119: out<=1;
   30120: out<=1;
   30121: out<=0;
   30122: out<=1;
   30123: out<=0;
   30124: out<=1;
   30125: out<=1;
   30126: out<=0;
   30127: out<=0;
   30128: out<=0;
   30129: out<=1;
   30130: out<=1;
   30131: out<=0;
   30132: out<=1;
   30133: out<=1;
   30134: out<=1;
   30135: out<=1;
   30136: out<=1;
   30137: out<=1;
   30138: out<=0;
   30139: out<=0;
   30140: out<=0;
   30141: out<=1;
   30142: out<=0;
   30143: out<=1;
   30144: out<=0;
   30145: out<=1;
   30146: out<=0;
   30147: out<=1;
   30148: out<=1;
   30149: out<=1;
   30150: out<=0;
   30151: out<=0;
   30152: out<=0;
   30153: out<=0;
   30154: out<=0;
   30155: out<=0;
   30156: out<=1;
   30157: out<=0;
   30158: out<=0;
   30159: out<=1;
   30160: out<=0;
   30161: out<=0;
   30162: out<=1;
   30163: out<=1;
   30164: out<=0;
   30165: out<=1;
   30166: out<=0;
   30167: out<=1;
   30168: out<=1;
   30169: out<=0;
   30170: out<=0;
   30171: out<=1;
   30172: out<=1;
   30173: out<=1;
   30174: out<=1;
   30175: out<=1;
   30176: out<=0;
   30177: out<=0;
   30178: out<=0;
   30179: out<=0;
   30180: out<=0;
   30181: out<=1;
   30182: out<=1;
   30183: out<=0;
   30184: out<=0;
   30185: out<=1;
   30186: out<=0;
   30187: out<=1;
   30188: out<=0;
   30189: out<=0;
   30190: out<=1;
   30191: out<=1;
   30192: out<=0;
   30193: out<=1;
   30194: out<=1;
   30195: out<=0;
   30196: out<=1;
   30197: out<=1;
   30198: out<=1;
   30199: out<=1;
   30200: out<=1;
   30201: out<=1;
   30202: out<=0;
   30203: out<=0;
   30204: out<=0;
   30205: out<=1;
   30206: out<=0;
   30207: out<=1;
   30208: out<=0;
   30209: out<=1;
   30210: out<=1;
   30211: out<=0;
   30212: out<=1;
   30213: out<=1;
   30214: out<=1;
   30215: out<=1;
   30216: out<=1;
   30217: out<=1;
   30218: out<=0;
   30219: out<=0;
   30220: out<=0;
   30221: out<=1;
   30222: out<=0;
   30223: out<=1;
   30224: out<=0;
   30225: out<=0;
   30226: out<=0;
   30227: out<=0;
   30228: out<=0;
   30229: out<=1;
   30230: out<=1;
   30231: out<=0;
   30232: out<=0;
   30233: out<=1;
   30234: out<=0;
   30235: out<=1;
   30236: out<=0;
   30237: out<=0;
   30238: out<=1;
   30239: out<=1;
   30240: out<=0;
   30241: out<=0;
   30242: out<=1;
   30243: out<=1;
   30244: out<=0;
   30245: out<=1;
   30246: out<=0;
   30247: out<=1;
   30248: out<=1;
   30249: out<=0;
   30250: out<=0;
   30251: out<=1;
   30252: out<=1;
   30253: out<=1;
   30254: out<=1;
   30255: out<=1;
   30256: out<=0;
   30257: out<=1;
   30258: out<=0;
   30259: out<=1;
   30260: out<=1;
   30261: out<=1;
   30262: out<=0;
   30263: out<=0;
   30264: out<=0;
   30265: out<=0;
   30266: out<=0;
   30267: out<=0;
   30268: out<=1;
   30269: out<=0;
   30270: out<=0;
   30271: out<=1;
   30272: out<=0;
   30273: out<=1;
   30274: out<=1;
   30275: out<=0;
   30276: out<=1;
   30277: out<=1;
   30278: out<=1;
   30279: out<=1;
   30280: out<=1;
   30281: out<=1;
   30282: out<=0;
   30283: out<=0;
   30284: out<=0;
   30285: out<=1;
   30286: out<=0;
   30287: out<=1;
   30288: out<=1;
   30289: out<=1;
   30290: out<=1;
   30291: out<=1;
   30292: out<=1;
   30293: out<=0;
   30294: out<=0;
   30295: out<=1;
   30296: out<=1;
   30297: out<=0;
   30298: out<=1;
   30299: out<=0;
   30300: out<=1;
   30301: out<=1;
   30302: out<=0;
   30303: out<=0;
   30304: out<=1;
   30305: out<=1;
   30306: out<=0;
   30307: out<=0;
   30308: out<=1;
   30309: out<=0;
   30310: out<=1;
   30311: out<=0;
   30312: out<=0;
   30313: out<=1;
   30314: out<=1;
   30315: out<=0;
   30316: out<=0;
   30317: out<=0;
   30318: out<=0;
   30319: out<=0;
   30320: out<=0;
   30321: out<=1;
   30322: out<=0;
   30323: out<=1;
   30324: out<=1;
   30325: out<=1;
   30326: out<=0;
   30327: out<=0;
   30328: out<=0;
   30329: out<=0;
   30330: out<=0;
   30331: out<=0;
   30332: out<=1;
   30333: out<=0;
   30334: out<=0;
   30335: out<=1;
   30336: out<=0;
   30337: out<=1;
   30338: out<=1;
   30339: out<=0;
   30340: out<=1;
   30341: out<=1;
   30342: out<=1;
   30343: out<=1;
   30344: out<=1;
   30345: out<=1;
   30346: out<=0;
   30347: out<=0;
   30348: out<=0;
   30349: out<=1;
   30350: out<=0;
   30351: out<=1;
   30352: out<=1;
   30353: out<=1;
   30354: out<=1;
   30355: out<=1;
   30356: out<=1;
   30357: out<=0;
   30358: out<=0;
   30359: out<=1;
   30360: out<=1;
   30361: out<=0;
   30362: out<=1;
   30363: out<=0;
   30364: out<=1;
   30365: out<=1;
   30366: out<=0;
   30367: out<=0;
   30368: out<=0;
   30369: out<=0;
   30370: out<=1;
   30371: out<=1;
   30372: out<=0;
   30373: out<=1;
   30374: out<=0;
   30375: out<=1;
   30376: out<=1;
   30377: out<=0;
   30378: out<=0;
   30379: out<=1;
   30380: out<=1;
   30381: out<=1;
   30382: out<=1;
   30383: out<=1;
   30384: out<=1;
   30385: out<=0;
   30386: out<=1;
   30387: out<=0;
   30388: out<=0;
   30389: out<=0;
   30390: out<=1;
   30391: out<=1;
   30392: out<=1;
   30393: out<=1;
   30394: out<=1;
   30395: out<=1;
   30396: out<=0;
   30397: out<=1;
   30398: out<=1;
   30399: out<=0;
   30400: out<=0;
   30401: out<=1;
   30402: out<=1;
   30403: out<=0;
   30404: out<=1;
   30405: out<=1;
   30406: out<=1;
   30407: out<=1;
   30408: out<=1;
   30409: out<=1;
   30410: out<=0;
   30411: out<=0;
   30412: out<=0;
   30413: out<=1;
   30414: out<=0;
   30415: out<=1;
   30416: out<=0;
   30417: out<=0;
   30418: out<=0;
   30419: out<=0;
   30420: out<=0;
   30421: out<=1;
   30422: out<=1;
   30423: out<=0;
   30424: out<=0;
   30425: out<=1;
   30426: out<=0;
   30427: out<=1;
   30428: out<=0;
   30429: out<=0;
   30430: out<=1;
   30431: out<=1;
   30432: out<=1;
   30433: out<=1;
   30434: out<=0;
   30435: out<=0;
   30436: out<=1;
   30437: out<=0;
   30438: out<=1;
   30439: out<=0;
   30440: out<=0;
   30441: out<=1;
   30442: out<=1;
   30443: out<=0;
   30444: out<=0;
   30445: out<=0;
   30446: out<=0;
   30447: out<=0;
   30448: out<=1;
   30449: out<=0;
   30450: out<=1;
   30451: out<=0;
   30452: out<=0;
   30453: out<=0;
   30454: out<=1;
   30455: out<=1;
   30456: out<=1;
   30457: out<=1;
   30458: out<=1;
   30459: out<=1;
   30460: out<=0;
   30461: out<=1;
   30462: out<=1;
   30463: out<=0;
   30464: out<=1;
   30465: out<=1;
   30466: out<=1;
   30467: out<=1;
   30468: out<=1;
   30469: out<=0;
   30470: out<=0;
   30471: out<=1;
   30472: out<=1;
   30473: out<=0;
   30474: out<=1;
   30475: out<=0;
   30476: out<=1;
   30477: out<=1;
   30478: out<=0;
   30479: out<=0;
   30480: out<=0;
   30481: out<=1;
   30482: out<=1;
   30483: out<=0;
   30484: out<=1;
   30485: out<=1;
   30486: out<=1;
   30487: out<=1;
   30488: out<=1;
   30489: out<=1;
   30490: out<=0;
   30491: out<=0;
   30492: out<=0;
   30493: out<=1;
   30494: out<=0;
   30495: out<=1;
   30496: out<=0;
   30497: out<=1;
   30498: out<=0;
   30499: out<=1;
   30500: out<=1;
   30501: out<=1;
   30502: out<=0;
   30503: out<=0;
   30504: out<=0;
   30505: out<=0;
   30506: out<=0;
   30507: out<=0;
   30508: out<=1;
   30509: out<=0;
   30510: out<=0;
   30511: out<=1;
   30512: out<=1;
   30513: out<=1;
   30514: out<=0;
   30515: out<=0;
   30516: out<=1;
   30517: out<=0;
   30518: out<=1;
   30519: out<=0;
   30520: out<=0;
   30521: out<=1;
   30522: out<=1;
   30523: out<=0;
   30524: out<=0;
   30525: out<=0;
   30526: out<=0;
   30527: out<=0;
   30528: out<=0;
   30529: out<=0;
   30530: out<=0;
   30531: out<=0;
   30532: out<=0;
   30533: out<=1;
   30534: out<=1;
   30535: out<=0;
   30536: out<=0;
   30537: out<=1;
   30538: out<=0;
   30539: out<=1;
   30540: out<=0;
   30541: out<=0;
   30542: out<=1;
   30543: out<=1;
   30544: out<=0;
   30545: out<=1;
   30546: out<=1;
   30547: out<=0;
   30548: out<=1;
   30549: out<=1;
   30550: out<=1;
   30551: out<=1;
   30552: out<=1;
   30553: out<=1;
   30554: out<=0;
   30555: out<=0;
   30556: out<=0;
   30557: out<=1;
   30558: out<=0;
   30559: out<=1;
   30560: out<=0;
   30561: out<=1;
   30562: out<=0;
   30563: out<=1;
   30564: out<=1;
   30565: out<=1;
   30566: out<=0;
   30567: out<=0;
   30568: out<=0;
   30569: out<=0;
   30570: out<=0;
   30571: out<=0;
   30572: out<=1;
   30573: out<=0;
   30574: out<=0;
   30575: out<=1;
   30576: out<=0;
   30577: out<=0;
   30578: out<=1;
   30579: out<=1;
   30580: out<=0;
   30581: out<=1;
   30582: out<=0;
   30583: out<=1;
   30584: out<=1;
   30585: out<=0;
   30586: out<=0;
   30587: out<=1;
   30588: out<=1;
   30589: out<=1;
   30590: out<=1;
   30591: out<=1;
   30592: out<=0;
   30593: out<=0;
   30594: out<=0;
   30595: out<=0;
   30596: out<=0;
   30597: out<=1;
   30598: out<=1;
   30599: out<=0;
   30600: out<=0;
   30601: out<=1;
   30602: out<=0;
   30603: out<=1;
   30604: out<=0;
   30605: out<=0;
   30606: out<=1;
   30607: out<=1;
   30608: out<=0;
   30609: out<=1;
   30610: out<=1;
   30611: out<=0;
   30612: out<=1;
   30613: out<=1;
   30614: out<=1;
   30615: out<=1;
   30616: out<=1;
   30617: out<=1;
   30618: out<=0;
   30619: out<=0;
   30620: out<=0;
   30621: out<=1;
   30622: out<=0;
   30623: out<=1;
   30624: out<=1;
   30625: out<=0;
   30626: out<=1;
   30627: out<=0;
   30628: out<=0;
   30629: out<=0;
   30630: out<=1;
   30631: out<=1;
   30632: out<=1;
   30633: out<=1;
   30634: out<=1;
   30635: out<=1;
   30636: out<=0;
   30637: out<=1;
   30638: out<=1;
   30639: out<=0;
   30640: out<=1;
   30641: out<=1;
   30642: out<=0;
   30643: out<=0;
   30644: out<=1;
   30645: out<=0;
   30646: out<=1;
   30647: out<=0;
   30648: out<=0;
   30649: out<=1;
   30650: out<=1;
   30651: out<=0;
   30652: out<=0;
   30653: out<=0;
   30654: out<=0;
   30655: out<=0;
   30656: out<=1;
   30657: out<=1;
   30658: out<=1;
   30659: out<=1;
   30660: out<=1;
   30661: out<=0;
   30662: out<=0;
   30663: out<=1;
   30664: out<=1;
   30665: out<=0;
   30666: out<=1;
   30667: out<=0;
   30668: out<=1;
   30669: out<=1;
   30670: out<=0;
   30671: out<=0;
   30672: out<=0;
   30673: out<=1;
   30674: out<=1;
   30675: out<=0;
   30676: out<=1;
   30677: out<=1;
   30678: out<=1;
   30679: out<=1;
   30680: out<=1;
   30681: out<=1;
   30682: out<=0;
   30683: out<=0;
   30684: out<=0;
   30685: out<=1;
   30686: out<=0;
   30687: out<=1;
   30688: out<=1;
   30689: out<=0;
   30690: out<=1;
   30691: out<=0;
   30692: out<=0;
   30693: out<=0;
   30694: out<=1;
   30695: out<=1;
   30696: out<=1;
   30697: out<=1;
   30698: out<=1;
   30699: out<=1;
   30700: out<=0;
   30701: out<=1;
   30702: out<=1;
   30703: out<=0;
   30704: out<=0;
   30705: out<=0;
   30706: out<=1;
   30707: out<=1;
   30708: out<=0;
   30709: out<=1;
   30710: out<=0;
   30711: out<=1;
   30712: out<=1;
   30713: out<=0;
   30714: out<=0;
   30715: out<=1;
   30716: out<=1;
   30717: out<=1;
   30718: out<=1;
   30719: out<=1;
   30720: out<=1;
   30721: out<=1;
   30722: out<=1;
   30723: out<=1;
   30724: out<=1;
   30725: out<=0;
   30726: out<=0;
   30727: out<=1;
   30728: out<=0;
   30729: out<=1;
   30730: out<=0;
   30731: out<=1;
   30732: out<=0;
   30733: out<=0;
   30734: out<=1;
   30735: out<=1;
   30736: out<=0;
   30737: out<=1;
   30738: out<=1;
   30739: out<=0;
   30740: out<=1;
   30741: out<=1;
   30742: out<=1;
   30743: out<=1;
   30744: out<=0;
   30745: out<=0;
   30746: out<=1;
   30747: out<=1;
   30748: out<=1;
   30749: out<=0;
   30750: out<=1;
   30751: out<=0;
   30752: out<=1;
   30753: out<=0;
   30754: out<=1;
   30755: out<=0;
   30756: out<=0;
   30757: out<=0;
   30758: out<=1;
   30759: out<=1;
   30760: out<=0;
   30761: out<=0;
   30762: out<=0;
   30763: out<=0;
   30764: out<=1;
   30765: out<=0;
   30766: out<=0;
   30767: out<=1;
   30768: out<=0;
   30769: out<=0;
   30770: out<=1;
   30771: out<=1;
   30772: out<=0;
   30773: out<=1;
   30774: out<=0;
   30775: out<=1;
   30776: out<=0;
   30777: out<=1;
   30778: out<=1;
   30779: out<=0;
   30780: out<=0;
   30781: out<=0;
   30782: out<=0;
   30783: out<=0;
   30784: out<=0;
   30785: out<=0;
   30786: out<=0;
   30787: out<=0;
   30788: out<=0;
   30789: out<=1;
   30790: out<=1;
   30791: out<=0;
   30792: out<=1;
   30793: out<=0;
   30794: out<=1;
   30795: out<=0;
   30796: out<=1;
   30797: out<=1;
   30798: out<=0;
   30799: out<=0;
   30800: out<=0;
   30801: out<=1;
   30802: out<=1;
   30803: out<=0;
   30804: out<=1;
   30805: out<=1;
   30806: out<=1;
   30807: out<=1;
   30808: out<=0;
   30809: out<=0;
   30810: out<=1;
   30811: out<=1;
   30812: out<=1;
   30813: out<=0;
   30814: out<=1;
   30815: out<=0;
   30816: out<=1;
   30817: out<=0;
   30818: out<=1;
   30819: out<=0;
   30820: out<=0;
   30821: out<=0;
   30822: out<=1;
   30823: out<=1;
   30824: out<=0;
   30825: out<=0;
   30826: out<=0;
   30827: out<=0;
   30828: out<=1;
   30829: out<=0;
   30830: out<=0;
   30831: out<=1;
   30832: out<=1;
   30833: out<=1;
   30834: out<=0;
   30835: out<=0;
   30836: out<=1;
   30837: out<=0;
   30838: out<=1;
   30839: out<=0;
   30840: out<=1;
   30841: out<=0;
   30842: out<=0;
   30843: out<=1;
   30844: out<=1;
   30845: out<=1;
   30846: out<=1;
   30847: out<=1;
   30848: out<=0;
   30849: out<=0;
   30850: out<=0;
   30851: out<=0;
   30852: out<=0;
   30853: out<=1;
   30854: out<=1;
   30855: out<=0;
   30856: out<=1;
   30857: out<=0;
   30858: out<=1;
   30859: out<=0;
   30860: out<=1;
   30861: out<=1;
   30862: out<=0;
   30863: out<=0;
   30864: out<=0;
   30865: out<=1;
   30866: out<=1;
   30867: out<=0;
   30868: out<=1;
   30869: out<=1;
   30870: out<=1;
   30871: out<=1;
   30872: out<=0;
   30873: out<=0;
   30874: out<=1;
   30875: out<=1;
   30876: out<=1;
   30877: out<=0;
   30878: out<=1;
   30879: out<=0;
   30880: out<=0;
   30881: out<=1;
   30882: out<=0;
   30883: out<=1;
   30884: out<=1;
   30885: out<=1;
   30886: out<=0;
   30887: out<=0;
   30888: out<=1;
   30889: out<=1;
   30890: out<=1;
   30891: out<=1;
   30892: out<=0;
   30893: out<=1;
   30894: out<=1;
   30895: out<=0;
   30896: out<=0;
   30897: out<=0;
   30898: out<=1;
   30899: out<=1;
   30900: out<=0;
   30901: out<=1;
   30902: out<=0;
   30903: out<=1;
   30904: out<=0;
   30905: out<=1;
   30906: out<=1;
   30907: out<=0;
   30908: out<=0;
   30909: out<=0;
   30910: out<=0;
   30911: out<=0;
   30912: out<=1;
   30913: out<=1;
   30914: out<=1;
   30915: out<=1;
   30916: out<=1;
   30917: out<=0;
   30918: out<=0;
   30919: out<=1;
   30920: out<=0;
   30921: out<=1;
   30922: out<=0;
   30923: out<=1;
   30924: out<=0;
   30925: out<=0;
   30926: out<=1;
   30927: out<=1;
   30928: out<=0;
   30929: out<=1;
   30930: out<=1;
   30931: out<=0;
   30932: out<=1;
   30933: out<=1;
   30934: out<=1;
   30935: out<=1;
   30936: out<=0;
   30937: out<=0;
   30938: out<=1;
   30939: out<=1;
   30940: out<=1;
   30941: out<=0;
   30942: out<=1;
   30943: out<=0;
   30944: out<=0;
   30945: out<=1;
   30946: out<=0;
   30947: out<=1;
   30948: out<=1;
   30949: out<=1;
   30950: out<=0;
   30951: out<=0;
   30952: out<=1;
   30953: out<=1;
   30954: out<=1;
   30955: out<=1;
   30956: out<=0;
   30957: out<=1;
   30958: out<=1;
   30959: out<=0;
   30960: out<=1;
   30961: out<=1;
   30962: out<=0;
   30963: out<=0;
   30964: out<=1;
   30965: out<=0;
   30966: out<=1;
   30967: out<=0;
   30968: out<=1;
   30969: out<=0;
   30970: out<=0;
   30971: out<=1;
   30972: out<=1;
   30973: out<=1;
   30974: out<=1;
   30975: out<=1;
   30976: out<=0;
   30977: out<=1;
   30978: out<=1;
   30979: out<=0;
   30980: out<=1;
   30981: out<=1;
   30982: out<=1;
   30983: out<=1;
   30984: out<=0;
   30985: out<=0;
   30986: out<=1;
   30987: out<=1;
   30988: out<=1;
   30989: out<=0;
   30990: out<=1;
   30991: out<=0;
   30992: out<=0;
   30993: out<=0;
   30994: out<=0;
   30995: out<=0;
   30996: out<=0;
   30997: out<=1;
   30998: out<=1;
   30999: out<=0;
   31000: out<=1;
   31001: out<=0;
   31002: out<=1;
   31003: out<=0;
   31004: out<=1;
   31005: out<=1;
   31006: out<=0;
   31007: out<=0;
   31008: out<=1;
   31009: out<=1;
   31010: out<=0;
   31011: out<=0;
   31012: out<=1;
   31013: out<=0;
   31014: out<=1;
   31015: out<=0;
   31016: out<=1;
   31017: out<=0;
   31018: out<=0;
   31019: out<=1;
   31020: out<=1;
   31021: out<=1;
   31022: out<=1;
   31023: out<=1;
   31024: out<=1;
   31025: out<=0;
   31026: out<=1;
   31027: out<=0;
   31028: out<=0;
   31029: out<=0;
   31030: out<=1;
   31031: out<=1;
   31032: out<=0;
   31033: out<=0;
   31034: out<=0;
   31035: out<=0;
   31036: out<=1;
   31037: out<=0;
   31038: out<=0;
   31039: out<=1;
   31040: out<=0;
   31041: out<=1;
   31042: out<=1;
   31043: out<=0;
   31044: out<=1;
   31045: out<=1;
   31046: out<=1;
   31047: out<=1;
   31048: out<=0;
   31049: out<=0;
   31050: out<=1;
   31051: out<=1;
   31052: out<=1;
   31053: out<=0;
   31054: out<=1;
   31055: out<=0;
   31056: out<=1;
   31057: out<=1;
   31058: out<=1;
   31059: out<=1;
   31060: out<=1;
   31061: out<=0;
   31062: out<=0;
   31063: out<=1;
   31064: out<=0;
   31065: out<=1;
   31066: out<=0;
   31067: out<=1;
   31068: out<=0;
   31069: out<=0;
   31070: out<=1;
   31071: out<=1;
   31072: out<=0;
   31073: out<=0;
   31074: out<=1;
   31075: out<=1;
   31076: out<=0;
   31077: out<=1;
   31078: out<=0;
   31079: out<=1;
   31080: out<=0;
   31081: out<=1;
   31082: out<=1;
   31083: out<=0;
   31084: out<=0;
   31085: out<=0;
   31086: out<=0;
   31087: out<=0;
   31088: out<=1;
   31089: out<=0;
   31090: out<=1;
   31091: out<=0;
   31092: out<=0;
   31093: out<=0;
   31094: out<=1;
   31095: out<=1;
   31096: out<=0;
   31097: out<=0;
   31098: out<=0;
   31099: out<=0;
   31100: out<=1;
   31101: out<=0;
   31102: out<=0;
   31103: out<=1;
   31104: out<=0;
   31105: out<=1;
   31106: out<=1;
   31107: out<=0;
   31108: out<=1;
   31109: out<=1;
   31110: out<=1;
   31111: out<=1;
   31112: out<=0;
   31113: out<=0;
   31114: out<=1;
   31115: out<=1;
   31116: out<=1;
   31117: out<=0;
   31118: out<=1;
   31119: out<=0;
   31120: out<=1;
   31121: out<=1;
   31122: out<=1;
   31123: out<=1;
   31124: out<=1;
   31125: out<=0;
   31126: out<=0;
   31127: out<=1;
   31128: out<=0;
   31129: out<=1;
   31130: out<=0;
   31131: out<=1;
   31132: out<=0;
   31133: out<=0;
   31134: out<=1;
   31135: out<=1;
   31136: out<=1;
   31137: out<=1;
   31138: out<=0;
   31139: out<=0;
   31140: out<=1;
   31141: out<=0;
   31142: out<=1;
   31143: out<=0;
   31144: out<=1;
   31145: out<=0;
   31146: out<=0;
   31147: out<=1;
   31148: out<=1;
   31149: out<=1;
   31150: out<=1;
   31151: out<=1;
   31152: out<=0;
   31153: out<=1;
   31154: out<=0;
   31155: out<=1;
   31156: out<=1;
   31157: out<=1;
   31158: out<=0;
   31159: out<=0;
   31160: out<=1;
   31161: out<=1;
   31162: out<=1;
   31163: out<=1;
   31164: out<=0;
   31165: out<=1;
   31166: out<=1;
   31167: out<=0;
   31168: out<=0;
   31169: out<=1;
   31170: out<=1;
   31171: out<=0;
   31172: out<=1;
   31173: out<=1;
   31174: out<=1;
   31175: out<=1;
   31176: out<=0;
   31177: out<=0;
   31178: out<=1;
   31179: out<=1;
   31180: out<=1;
   31181: out<=0;
   31182: out<=1;
   31183: out<=0;
   31184: out<=0;
   31185: out<=0;
   31186: out<=0;
   31187: out<=0;
   31188: out<=0;
   31189: out<=1;
   31190: out<=1;
   31191: out<=0;
   31192: out<=1;
   31193: out<=0;
   31194: out<=1;
   31195: out<=0;
   31196: out<=1;
   31197: out<=1;
   31198: out<=0;
   31199: out<=0;
   31200: out<=0;
   31201: out<=0;
   31202: out<=1;
   31203: out<=1;
   31204: out<=0;
   31205: out<=1;
   31206: out<=0;
   31207: out<=1;
   31208: out<=0;
   31209: out<=1;
   31210: out<=1;
   31211: out<=0;
   31212: out<=0;
   31213: out<=0;
   31214: out<=0;
   31215: out<=0;
   31216: out<=0;
   31217: out<=1;
   31218: out<=0;
   31219: out<=1;
   31220: out<=1;
   31221: out<=1;
   31222: out<=0;
   31223: out<=0;
   31224: out<=1;
   31225: out<=1;
   31226: out<=1;
   31227: out<=1;
   31228: out<=0;
   31229: out<=1;
   31230: out<=1;
   31231: out<=0;
   31232: out<=0;
   31233: out<=1;
   31234: out<=0;
   31235: out<=1;
   31236: out<=1;
   31237: out<=1;
   31238: out<=0;
   31239: out<=0;
   31240: out<=1;
   31241: out<=1;
   31242: out<=1;
   31243: out<=1;
   31244: out<=0;
   31245: out<=1;
   31246: out<=1;
   31247: out<=0;
   31248: out<=0;
   31249: out<=0;
   31250: out<=1;
   31251: out<=1;
   31252: out<=0;
   31253: out<=1;
   31254: out<=0;
   31255: out<=1;
   31256: out<=0;
   31257: out<=1;
   31258: out<=1;
   31259: out<=0;
   31260: out<=0;
   31261: out<=0;
   31262: out<=0;
   31263: out<=0;
   31264: out<=0;
   31265: out<=0;
   31266: out<=0;
   31267: out<=0;
   31268: out<=0;
   31269: out<=1;
   31270: out<=1;
   31271: out<=0;
   31272: out<=1;
   31273: out<=0;
   31274: out<=1;
   31275: out<=0;
   31276: out<=1;
   31277: out<=1;
   31278: out<=0;
   31279: out<=0;
   31280: out<=0;
   31281: out<=1;
   31282: out<=1;
   31283: out<=0;
   31284: out<=1;
   31285: out<=1;
   31286: out<=1;
   31287: out<=1;
   31288: out<=0;
   31289: out<=0;
   31290: out<=1;
   31291: out<=1;
   31292: out<=1;
   31293: out<=0;
   31294: out<=1;
   31295: out<=0;
   31296: out<=0;
   31297: out<=1;
   31298: out<=0;
   31299: out<=1;
   31300: out<=1;
   31301: out<=1;
   31302: out<=0;
   31303: out<=0;
   31304: out<=1;
   31305: out<=1;
   31306: out<=1;
   31307: out<=1;
   31308: out<=0;
   31309: out<=1;
   31310: out<=1;
   31311: out<=0;
   31312: out<=1;
   31313: out<=1;
   31314: out<=0;
   31315: out<=0;
   31316: out<=1;
   31317: out<=0;
   31318: out<=1;
   31319: out<=0;
   31320: out<=1;
   31321: out<=0;
   31322: out<=0;
   31323: out<=1;
   31324: out<=1;
   31325: out<=1;
   31326: out<=1;
   31327: out<=1;
   31328: out<=1;
   31329: out<=1;
   31330: out<=1;
   31331: out<=1;
   31332: out<=1;
   31333: out<=0;
   31334: out<=0;
   31335: out<=1;
   31336: out<=0;
   31337: out<=1;
   31338: out<=0;
   31339: out<=1;
   31340: out<=0;
   31341: out<=0;
   31342: out<=1;
   31343: out<=1;
   31344: out<=0;
   31345: out<=1;
   31346: out<=1;
   31347: out<=0;
   31348: out<=1;
   31349: out<=1;
   31350: out<=1;
   31351: out<=1;
   31352: out<=0;
   31353: out<=0;
   31354: out<=1;
   31355: out<=1;
   31356: out<=1;
   31357: out<=0;
   31358: out<=1;
   31359: out<=0;
   31360: out<=1;
   31361: out<=0;
   31362: out<=1;
   31363: out<=0;
   31364: out<=0;
   31365: out<=0;
   31366: out<=1;
   31367: out<=1;
   31368: out<=0;
   31369: out<=0;
   31370: out<=0;
   31371: out<=0;
   31372: out<=1;
   31373: out<=0;
   31374: out<=0;
   31375: out<=1;
   31376: out<=0;
   31377: out<=0;
   31378: out<=1;
   31379: out<=1;
   31380: out<=0;
   31381: out<=1;
   31382: out<=0;
   31383: out<=1;
   31384: out<=0;
   31385: out<=1;
   31386: out<=1;
   31387: out<=0;
   31388: out<=0;
   31389: out<=0;
   31390: out<=0;
   31391: out<=0;
   31392: out<=1;
   31393: out<=1;
   31394: out<=1;
   31395: out<=1;
   31396: out<=1;
   31397: out<=0;
   31398: out<=0;
   31399: out<=1;
   31400: out<=0;
   31401: out<=1;
   31402: out<=0;
   31403: out<=1;
   31404: out<=0;
   31405: out<=0;
   31406: out<=1;
   31407: out<=1;
   31408: out<=0;
   31409: out<=1;
   31410: out<=1;
   31411: out<=0;
   31412: out<=1;
   31413: out<=1;
   31414: out<=1;
   31415: out<=1;
   31416: out<=0;
   31417: out<=0;
   31418: out<=1;
   31419: out<=1;
   31420: out<=1;
   31421: out<=0;
   31422: out<=1;
   31423: out<=0;
   31424: out<=1;
   31425: out<=0;
   31426: out<=1;
   31427: out<=0;
   31428: out<=0;
   31429: out<=0;
   31430: out<=1;
   31431: out<=1;
   31432: out<=0;
   31433: out<=0;
   31434: out<=0;
   31435: out<=0;
   31436: out<=1;
   31437: out<=0;
   31438: out<=0;
   31439: out<=1;
   31440: out<=1;
   31441: out<=1;
   31442: out<=0;
   31443: out<=0;
   31444: out<=1;
   31445: out<=0;
   31446: out<=1;
   31447: out<=0;
   31448: out<=1;
   31449: out<=0;
   31450: out<=0;
   31451: out<=1;
   31452: out<=1;
   31453: out<=1;
   31454: out<=1;
   31455: out<=1;
   31456: out<=0;
   31457: out<=0;
   31458: out<=0;
   31459: out<=0;
   31460: out<=0;
   31461: out<=1;
   31462: out<=1;
   31463: out<=0;
   31464: out<=1;
   31465: out<=0;
   31466: out<=1;
   31467: out<=0;
   31468: out<=1;
   31469: out<=1;
   31470: out<=0;
   31471: out<=0;
   31472: out<=0;
   31473: out<=1;
   31474: out<=1;
   31475: out<=0;
   31476: out<=1;
   31477: out<=1;
   31478: out<=1;
   31479: out<=1;
   31480: out<=0;
   31481: out<=0;
   31482: out<=1;
   31483: out<=1;
   31484: out<=1;
   31485: out<=0;
   31486: out<=1;
   31487: out<=0;
   31488: out<=1;
   31489: out<=1;
   31490: out<=0;
   31491: out<=0;
   31492: out<=1;
   31493: out<=0;
   31494: out<=1;
   31495: out<=0;
   31496: out<=1;
   31497: out<=0;
   31498: out<=0;
   31499: out<=1;
   31500: out<=1;
   31501: out<=1;
   31502: out<=1;
   31503: out<=1;
   31504: out<=0;
   31505: out<=1;
   31506: out<=0;
   31507: out<=1;
   31508: out<=1;
   31509: out<=1;
   31510: out<=0;
   31511: out<=0;
   31512: out<=1;
   31513: out<=1;
   31514: out<=1;
   31515: out<=1;
   31516: out<=0;
   31517: out<=1;
   31518: out<=1;
   31519: out<=0;
   31520: out<=0;
   31521: out<=1;
   31522: out<=1;
   31523: out<=0;
   31524: out<=1;
   31525: out<=1;
   31526: out<=1;
   31527: out<=1;
   31528: out<=0;
   31529: out<=0;
   31530: out<=1;
   31531: out<=1;
   31532: out<=1;
   31533: out<=0;
   31534: out<=1;
   31535: out<=0;
   31536: out<=1;
   31537: out<=1;
   31538: out<=1;
   31539: out<=1;
   31540: out<=1;
   31541: out<=0;
   31542: out<=0;
   31543: out<=1;
   31544: out<=0;
   31545: out<=1;
   31546: out<=0;
   31547: out<=1;
   31548: out<=0;
   31549: out<=0;
   31550: out<=1;
   31551: out<=1;
   31552: out<=0;
   31553: out<=0;
   31554: out<=1;
   31555: out<=1;
   31556: out<=0;
   31557: out<=1;
   31558: out<=0;
   31559: out<=1;
   31560: out<=0;
   31561: out<=1;
   31562: out<=1;
   31563: out<=0;
   31564: out<=0;
   31565: out<=0;
   31566: out<=0;
   31567: out<=0;
   31568: out<=0;
   31569: out<=1;
   31570: out<=0;
   31571: out<=1;
   31572: out<=1;
   31573: out<=1;
   31574: out<=0;
   31575: out<=0;
   31576: out<=1;
   31577: out<=1;
   31578: out<=1;
   31579: out<=1;
   31580: out<=0;
   31581: out<=1;
   31582: out<=1;
   31583: out<=0;
   31584: out<=0;
   31585: out<=1;
   31586: out<=1;
   31587: out<=0;
   31588: out<=1;
   31589: out<=1;
   31590: out<=1;
   31591: out<=1;
   31592: out<=0;
   31593: out<=0;
   31594: out<=1;
   31595: out<=1;
   31596: out<=1;
   31597: out<=0;
   31598: out<=1;
   31599: out<=0;
   31600: out<=0;
   31601: out<=0;
   31602: out<=0;
   31603: out<=0;
   31604: out<=0;
   31605: out<=1;
   31606: out<=1;
   31607: out<=0;
   31608: out<=1;
   31609: out<=0;
   31610: out<=1;
   31611: out<=0;
   31612: out<=1;
   31613: out<=1;
   31614: out<=0;
   31615: out<=0;
   31616: out<=1;
   31617: out<=1;
   31618: out<=0;
   31619: out<=0;
   31620: out<=1;
   31621: out<=0;
   31622: out<=1;
   31623: out<=0;
   31624: out<=1;
   31625: out<=0;
   31626: out<=0;
   31627: out<=1;
   31628: out<=1;
   31629: out<=1;
   31630: out<=1;
   31631: out<=1;
   31632: out<=1;
   31633: out<=0;
   31634: out<=1;
   31635: out<=0;
   31636: out<=0;
   31637: out<=0;
   31638: out<=1;
   31639: out<=1;
   31640: out<=0;
   31641: out<=0;
   31642: out<=0;
   31643: out<=0;
   31644: out<=1;
   31645: out<=0;
   31646: out<=0;
   31647: out<=1;
   31648: out<=0;
   31649: out<=1;
   31650: out<=1;
   31651: out<=0;
   31652: out<=1;
   31653: out<=1;
   31654: out<=1;
   31655: out<=1;
   31656: out<=0;
   31657: out<=0;
   31658: out<=1;
   31659: out<=1;
   31660: out<=1;
   31661: out<=0;
   31662: out<=1;
   31663: out<=0;
   31664: out<=0;
   31665: out<=0;
   31666: out<=0;
   31667: out<=0;
   31668: out<=0;
   31669: out<=1;
   31670: out<=1;
   31671: out<=0;
   31672: out<=1;
   31673: out<=0;
   31674: out<=1;
   31675: out<=0;
   31676: out<=1;
   31677: out<=1;
   31678: out<=0;
   31679: out<=0;
   31680: out<=0;
   31681: out<=0;
   31682: out<=1;
   31683: out<=1;
   31684: out<=0;
   31685: out<=1;
   31686: out<=0;
   31687: out<=1;
   31688: out<=0;
   31689: out<=1;
   31690: out<=1;
   31691: out<=0;
   31692: out<=0;
   31693: out<=0;
   31694: out<=0;
   31695: out<=0;
   31696: out<=1;
   31697: out<=0;
   31698: out<=1;
   31699: out<=0;
   31700: out<=0;
   31701: out<=0;
   31702: out<=1;
   31703: out<=1;
   31704: out<=0;
   31705: out<=0;
   31706: out<=0;
   31707: out<=0;
   31708: out<=1;
   31709: out<=0;
   31710: out<=0;
   31711: out<=1;
   31712: out<=0;
   31713: out<=1;
   31714: out<=1;
   31715: out<=0;
   31716: out<=1;
   31717: out<=1;
   31718: out<=1;
   31719: out<=1;
   31720: out<=0;
   31721: out<=0;
   31722: out<=1;
   31723: out<=1;
   31724: out<=1;
   31725: out<=0;
   31726: out<=1;
   31727: out<=0;
   31728: out<=1;
   31729: out<=1;
   31730: out<=1;
   31731: out<=1;
   31732: out<=1;
   31733: out<=0;
   31734: out<=0;
   31735: out<=1;
   31736: out<=0;
   31737: out<=1;
   31738: out<=0;
   31739: out<=1;
   31740: out<=0;
   31741: out<=0;
   31742: out<=1;
   31743: out<=1;
   31744: out<=1;
   31745: out<=0;
   31746: out<=0;
   31747: out<=1;
   31748: out<=1;
   31749: out<=1;
   31750: out<=1;
   31751: out<=1;
   31752: out<=0;
   31753: out<=0;
   31754: out<=1;
   31755: out<=1;
   31756: out<=0;
   31757: out<=1;
   31758: out<=0;
   31759: out<=1;
   31760: out<=0;
   31761: out<=0;
   31762: out<=0;
   31763: out<=0;
   31764: out<=1;
   31765: out<=0;
   31766: out<=0;
   31767: out<=1;
   31768: out<=0;
   31769: out<=1;
   31770: out<=0;
   31771: out<=1;
   31772: out<=1;
   31773: out<=1;
   31774: out<=0;
   31775: out<=0;
   31776: out<=1;
   31777: out<=1;
   31778: out<=0;
   31779: out<=0;
   31780: out<=0;
   31781: out<=1;
   31782: out<=0;
   31783: out<=1;
   31784: out<=0;
   31785: out<=1;
   31786: out<=1;
   31787: out<=0;
   31788: out<=1;
   31789: out<=1;
   31790: out<=1;
   31791: out<=1;
   31792: out<=0;
   31793: out<=1;
   31794: out<=0;
   31795: out<=1;
   31796: out<=0;
   31797: out<=0;
   31798: out<=1;
   31799: out<=1;
   31800: out<=0;
   31801: out<=0;
   31802: out<=0;
   31803: out<=0;
   31804: out<=0;
   31805: out<=1;
   31806: out<=1;
   31807: out<=0;
   31808: out<=1;
   31809: out<=0;
   31810: out<=0;
   31811: out<=1;
   31812: out<=1;
   31813: out<=1;
   31814: out<=1;
   31815: out<=1;
   31816: out<=0;
   31817: out<=0;
   31818: out<=1;
   31819: out<=1;
   31820: out<=0;
   31821: out<=1;
   31822: out<=0;
   31823: out<=1;
   31824: out<=1;
   31825: out<=1;
   31826: out<=1;
   31827: out<=1;
   31828: out<=0;
   31829: out<=1;
   31830: out<=1;
   31831: out<=0;
   31832: out<=1;
   31833: out<=0;
   31834: out<=1;
   31835: out<=0;
   31836: out<=0;
   31837: out<=0;
   31838: out<=1;
   31839: out<=1;
   31840: out<=0;
   31841: out<=0;
   31842: out<=1;
   31843: out<=1;
   31844: out<=1;
   31845: out<=0;
   31846: out<=1;
   31847: out<=0;
   31848: out<=1;
   31849: out<=0;
   31850: out<=0;
   31851: out<=1;
   31852: out<=0;
   31853: out<=0;
   31854: out<=0;
   31855: out<=0;
   31856: out<=0;
   31857: out<=1;
   31858: out<=0;
   31859: out<=1;
   31860: out<=0;
   31861: out<=0;
   31862: out<=1;
   31863: out<=1;
   31864: out<=0;
   31865: out<=0;
   31866: out<=0;
   31867: out<=0;
   31868: out<=0;
   31869: out<=1;
   31870: out<=1;
   31871: out<=0;
   31872: out<=1;
   31873: out<=0;
   31874: out<=0;
   31875: out<=1;
   31876: out<=1;
   31877: out<=1;
   31878: out<=1;
   31879: out<=1;
   31880: out<=0;
   31881: out<=0;
   31882: out<=1;
   31883: out<=1;
   31884: out<=0;
   31885: out<=1;
   31886: out<=0;
   31887: out<=1;
   31888: out<=1;
   31889: out<=1;
   31890: out<=1;
   31891: out<=1;
   31892: out<=0;
   31893: out<=1;
   31894: out<=1;
   31895: out<=0;
   31896: out<=1;
   31897: out<=0;
   31898: out<=1;
   31899: out<=0;
   31900: out<=0;
   31901: out<=0;
   31902: out<=1;
   31903: out<=1;
   31904: out<=1;
   31905: out<=1;
   31906: out<=0;
   31907: out<=0;
   31908: out<=0;
   31909: out<=1;
   31910: out<=0;
   31911: out<=1;
   31912: out<=0;
   31913: out<=1;
   31914: out<=1;
   31915: out<=0;
   31916: out<=1;
   31917: out<=1;
   31918: out<=1;
   31919: out<=1;
   31920: out<=1;
   31921: out<=0;
   31922: out<=1;
   31923: out<=0;
   31924: out<=1;
   31925: out<=1;
   31926: out<=0;
   31927: out<=0;
   31928: out<=1;
   31929: out<=1;
   31930: out<=1;
   31931: out<=1;
   31932: out<=1;
   31933: out<=0;
   31934: out<=0;
   31935: out<=1;
   31936: out<=1;
   31937: out<=0;
   31938: out<=0;
   31939: out<=1;
   31940: out<=1;
   31941: out<=1;
   31942: out<=1;
   31943: out<=1;
   31944: out<=0;
   31945: out<=0;
   31946: out<=1;
   31947: out<=1;
   31948: out<=0;
   31949: out<=1;
   31950: out<=0;
   31951: out<=1;
   31952: out<=0;
   31953: out<=0;
   31954: out<=0;
   31955: out<=0;
   31956: out<=1;
   31957: out<=0;
   31958: out<=0;
   31959: out<=1;
   31960: out<=0;
   31961: out<=1;
   31962: out<=0;
   31963: out<=1;
   31964: out<=1;
   31965: out<=1;
   31966: out<=0;
   31967: out<=0;
   31968: out<=0;
   31969: out<=0;
   31970: out<=1;
   31971: out<=1;
   31972: out<=1;
   31973: out<=0;
   31974: out<=1;
   31975: out<=0;
   31976: out<=1;
   31977: out<=0;
   31978: out<=0;
   31979: out<=1;
   31980: out<=0;
   31981: out<=0;
   31982: out<=0;
   31983: out<=0;
   31984: out<=1;
   31985: out<=0;
   31986: out<=1;
   31987: out<=0;
   31988: out<=1;
   31989: out<=1;
   31990: out<=0;
   31991: out<=0;
   31992: out<=1;
   31993: out<=1;
   31994: out<=1;
   31995: out<=1;
   31996: out<=1;
   31997: out<=0;
   31998: out<=0;
   31999: out<=1;
   32000: out<=1;
   32001: out<=1;
   32002: out<=1;
   32003: out<=1;
   32004: out<=0;
   32005: out<=1;
   32006: out<=1;
   32007: out<=0;
   32008: out<=1;
   32009: out<=0;
   32010: out<=1;
   32011: out<=0;
   32012: out<=0;
   32013: out<=0;
   32014: out<=1;
   32015: out<=1;
   32016: out<=1;
   32017: out<=0;
   32018: out<=0;
   32019: out<=1;
   32020: out<=1;
   32021: out<=1;
   32022: out<=1;
   32023: out<=1;
   32024: out<=0;
   32025: out<=0;
   32026: out<=1;
   32027: out<=1;
   32028: out<=0;
   32029: out<=1;
   32030: out<=0;
   32031: out<=1;
   32032: out<=0;
   32033: out<=1;
   32034: out<=0;
   32035: out<=1;
   32036: out<=0;
   32037: out<=0;
   32038: out<=1;
   32039: out<=1;
   32040: out<=0;
   32041: out<=0;
   32042: out<=0;
   32043: out<=0;
   32044: out<=0;
   32045: out<=1;
   32046: out<=1;
   32047: out<=0;
   32048: out<=0;
   32049: out<=0;
   32050: out<=1;
   32051: out<=1;
   32052: out<=1;
   32053: out<=0;
   32054: out<=1;
   32055: out<=0;
   32056: out<=1;
   32057: out<=0;
   32058: out<=0;
   32059: out<=1;
   32060: out<=0;
   32061: out<=0;
   32062: out<=0;
   32063: out<=0;
   32064: out<=0;
   32065: out<=0;
   32066: out<=0;
   32067: out<=0;
   32068: out<=1;
   32069: out<=0;
   32070: out<=0;
   32071: out<=1;
   32072: out<=0;
   32073: out<=1;
   32074: out<=0;
   32075: out<=1;
   32076: out<=1;
   32077: out<=1;
   32078: out<=0;
   32079: out<=0;
   32080: out<=1;
   32081: out<=0;
   32082: out<=0;
   32083: out<=1;
   32084: out<=1;
   32085: out<=1;
   32086: out<=1;
   32087: out<=1;
   32088: out<=0;
   32089: out<=0;
   32090: out<=1;
   32091: out<=1;
   32092: out<=0;
   32093: out<=1;
   32094: out<=0;
   32095: out<=1;
   32096: out<=0;
   32097: out<=1;
   32098: out<=0;
   32099: out<=1;
   32100: out<=0;
   32101: out<=0;
   32102: out<=1;
   32103: out<=1;
   32104: out<=0;
   32105: out<=0;
   32106: out<=0;
   32107: out<=0;
   32108: out<=0;
   32109: out<=1;
   32110: out<=1;
   32111: out<=0;
   32112: out<=1;
   32113: out<=1;
   32114: out<=0;
   32115: out<=0;
   32116: out<=0;
   32117: out<=1;
   32118: out<=0;
   32119: out<=1;
   32120: out<=0;
   32121: out<=1;
   32122: out<=1;
   32123: out<=0;
   32124: out<=1;
   32125: out<=1;
   32126: out<=1;
   32127: out<=1;
   32128: out<=0;
   32129: out<=0;
   32130: out<=0;
   32131: out<=0;
   32132: out<=1;
   32133: out<=0;
   32134: out<=0;
   32135: out<=1;
   32136: out<=0;
   32137: out<=1;
   32138: out<=0;
   32139: out<=1;
   32140: out<=1;
   32141: out<=1;
   32142: out<=0;
   32143: out<=0;
   32144: out<=1;
   32145: out<=0;
   32146: out<=0;
   32147: out<=1;
   32148: out<=1;
   32149: out<=1;
   32150: out<=1;
   32151: out<=1;
   32152: out<=0;
   32153: out<=0;
   32154: out<=1;
   32155: out<=1;
   32156: out<=0;
   32157: out<=1;
   32158: out<=0;
   32159: out<=1;
   32160: out<=1;
   32161: out<=0;
   32162: out<=1;
   32163: out<=0;
   32164: out<=1;
   32165: out<=1;
   32166: out<=0;
   32167: out<=0;
   32168: out<=1;
   32169: out<=1;
   32170: out<=1;
   32171: out<=1;
   32172: out<=1;
   32173: out<=0;
   32174: out<=0;
   32175: out<=1;
   32176: out<=0;
   32177: out<=0;
   32178: out<=1;
   32179: out<=1;
   32180: out<=1;
   32181: out<=0;
   32182: out<=1;
   32183: out<=0;
   32184: out<=1;
   32185: out<=0;
   32186: out<=0;
   32187: out<=1;
   32188: out<=0;
   32189: out<=0;
   32190: out<=0;
   32191: out<=0;
   32192: out<=1;
   32193: out<=1;
   32194: out<=1;
   32195: out<=1;
   32196: out<=0;
   32197: out<=1;
   32198: out<=1;
   32199: out<=0;
   32200: out<=1;
   32201: out<=0;
   32202: out<=1;
   32203: out<=0;
   32204: out<=0;
   32205: out<=0;
   32206: out<=1;
   32207: out<=1;
   32208: out<=1;
   32209: out<=0;
   32210: out<=0;
   32211: out<=1;
   32212: out<=1;
   32213: out<=1;
   32214: out<=1;
   32215: out<=1;
   32216: out<=0;
   32217: out<=0;
   32218: out<=1;
   32219: out<=1;
   32220: out<=0;
   32221: out<=1;
   32222: out<=0;
   32223: out<=1;
   32224: out<=1;
   32225: out<=0;
   32226: out<=1;
   32227: out<=0;
   32228: out<=1;
   32229: out<=1;
   32230: out<=0;
   32231: out<=0;
   32232: out<=1;
   32233: out<=1;
   32234: out<=1;
   32235: out<=1;
   32236: out<=1;
   32237: out<=0;
   32238: out<=0;
   32239: out<=1;
   32240: out<=1;
   32241: out<=1;
   32242: out<=0;
   32243: out<=0;
   32244: out<=0;
   32245: out<=1;
   32246: out<=0;
   32247: out<=1;
   32248: out<=0;
   32249: out<=1;
   32250: out<=1;
   32251: out<=0;
   32252: out<=1;
   32253: out<=1;
   32254: out<=1;
   32255: out<=1;
   32256: out<=1;
   32257: out<=1;
   32258: out<=0;
   32259: out<=0;
   32260: out<=0;
   32261: out<=1;
   32262: out<=0;
   32263: out<=1;
   32264: out<=0;
   32265: out<=1;
   32266: out<=1;
   32267: out<=0;
   32268: out<=1;
   32269: out<=1;
   32270: out<=1;
   32271: out<=1;
   32272: out<=1;
   32273: out<=0;
   32274: out<=1;
   32275: out<=0;
   32276: out<=1;
   32277: out<=1;
   32278: out<=0;
   32279: out<=0;
   32280: out<=1;
   32281: out<=1;
   32282: out<=1;
   32283: out<=1;
   32284: out<=1;
   32285: out<=0;
   32286: out<=0;
   32287: out<=1;
   32288: out<=1;
   32289: out<=0;
   32290: out<=0;
   32291: out<=1;
   32292: out<=1;
   32293: out<=1;
   32294: out<=1;
   32295: out<=1;
   32296: out<=0;
   32297: out<=0;
   32298: out<=1;
   32299: out<=1;
   32300: out<=0;
   32301: out<=1;
   32302: out<=0;
   32303: out<=1;
   32304: out<=1;
   32305: out<=1;
   32306: out<=1;
   32307: out<=1;
   32308: out<=0;
   32309: out<=1;
   32310: out<=1;
   32311: out<=0;
   32312: out<=1;
   32313: out<=0;
   32314: out<=1;
   32315: out<=0;
   32316: out<=0;
   32317: out<=0;
   32318: out<=1;
   32319: out<=1;
   32320: out<=0;
   32321: out<=0;
   32322: out<=1;
   32323: out<=1;
   32324: out<=1;
   32325: out<=0;
   32326: out<=1;
   32327: out<=0;
   32328: out<=1;
   32329: out<=0;
   32330: out<=0;
   32331: out<=1;
   32332: out<=0;
   32333: out<=0;
   32334: out<=0;
   32335: out<=0;
   32336: out<=1;
   32337: out<=0;
   32338: out<=1;
   32339: out<=0;
   32340: out<=1;
   32341: out<=1;
   32342: out<=0;
   32343: out<=0;
   32344: out<=1;
   32345: out<=1;
   32346: out<=1;
   32347: out<=1;
   32348: out<=1;
   32349: out<=0;
   32350: out<=0;
   32351: out<=1;
   32352: out<=1;
   32353: out<=0;
   32354: out<=0;
   32355: out<=1;
   32356: out<=1;
   32357: out<=1;
   32358: out<=1;
   32359: out<=1;
   32360: out<=0;
   32361: out<=0;
   32362: out<=1;
   32363: out<=1;
   32364: out<=0;
   32365: out<=1;
   32366: out<=0;
   32367: out<=1;
   32368: out<=0;
   32369: out<=0;
   32370: out<=0;
   32371: out<=0;
   32372: out<=1;
   32373: out<=0;
   32374: out<=0;
   32375: out<=1;
   32376: out<=0;
   32377: out<=1;
   32378: out<=0;
   32379: out<=1;
   32380: out<=1;
   32381: out<=1;
   32382: out<=0;
   32383: out<=0;
   32384: out<=1;
   32385: out<=1;
   32386: out<=0;
   32387: out<=0;
   32388: out<=0;
   32389: out<=1;
   32390: out<=0;
   32391: out<=1;
   32392: out<=0;
   32393: out<=1;
   32394: out<=1;
   32395: out<=0;
   32396: out<=1;
   32397: out<=1;
   32398: out<=1;
   32399: out<=1;
   32400: out<=0;
   32401: out<=1;
   32402: out<=0;
   32403: out<=1;
   32404: out<=0;
   32405: out<=0;
   32406: out<=1;
   32407: out<=1;
   32408: out<=0;
   32409: out<=0;
   32410: out<=0;
   32411: out<=0;
   32412: out<=0;
   32413: out<=1;
   32414: out<=1;
   32415: out<=0;
   32416: out<=1;
   32417: out<=0;
   32418: out<=0;
   32419: out<=1;
   32420: out<=1;
   32421: out<=1;
   32422: out<=1;
   32423: out<=1;
   32424: out<=0;
   32425: out<=0;
   32426: out<=1;
   32427: out<=1;
   32428: out<=0;
   32429: out<=1;
   32430: out<=0;
   32431: out<=1;
   32432: out<=0;
   32433: out<=0;
   32434: out<=0;
   32435: out<=0;
   32436: out<=1;
   32437: out<=0;
   32438: out<=0;
   32439: out<=1;
   32440: out<=0;
   32441: out<=1;
   32442: out<=0;
   32443: out<=1;
   32444: out<=1;
   32445: out<=1;
   32446: out<=0;
   32447: out<=0;
   32448: out<=0;
   32449: out<=0;
   32450: out<=1;
   32451: out<=1;
   32452: out<=1;
   32453: out<=0;
   32454: out<=1;
   32455: out<=0;
   32456: out<=1;
   32457: out<=0;
   32458: out<=0;
   32459: out<=1;
   32460: out<=0;
   32461: out<=0;
   32462: out<=0;
   32463: out<=0;
   32464: out<=0;
   32465: out<=1;
   32466: out<=0;
   32467: out<=1;
   32468: out<=0;
   32469: out<=0;
   32470: out<=1;
   32471: out<=1;
   32472: out<=0;
   32473: out<=0;
   32474: out<=0;
   32475: out<=0;
   32476: out<=0;
   32477: out<=1;
   32478: out<=1;
   32479: out<=0;
   32480: out<=1;
   32481: out<=0;
   32482: out<=0;
   32483: out<=1;
   32484: out<=1;
   32485: out<=1;
   32486: out<=1;
   32487: out<=1;
   32488: out<=0;
   32489: out<=0;
   32490: out<=1;
   32491: out<=1;
   32492: out<=0;
   32493: out<=1;
   32494: out<=0;
   32495: out<=1;
   32496: out<=1;
   32497: out<=1;
   32498: out<=1;
   32499: out<=1;
   32500: out<=0;
   32501: out<=1;
   32502: out<=1;
   32503: out<=0;
   32504: out<=1;
   32505: out<=0;
   32506: out<=1;
   32507: out<=0;
   32508: out<=0;
   32509: out<=0;
   32510: out<=1;
   32511: out<=1;
   32512: out<=1;
   32513: out<=0;
   32514: out<=1;
   32515: out<=0;
   32516: out<=1;
   32517: out<=1;
   32518: out<=0;
   32519: out<=0;
   32520: out<=1;
   32521: out<=1;
   32522: out<=1;
   32523: out<=1;
   32524: out<=1;
   32525: out<=0;
   32526: out<=0;
   32527: out<=1;
   32528: out<=0;
   32529: out<=0;
   32530: out<=1;
   32531: out<=1;
   32532: out<=1;
   32533: out<=0;
   32534: out<=1;
   32535: out<=0;
   32536: out<=1;
   32537: out<=0;
   32538: out<=0;
   32539: out<=1;
   32540: out<=0;
   32541: out<=0;
   32542: out<=0;
   32543: out<=0;
   32544: out<=0;
   32545: out<=0;
   32546: out<=0;
   32547: out<=0;
   32548: out<=1;
   32549: out<=0;
   32550: out<=0;
   32551: out<=1;
   32552: out<=0;
   32553: out<=1;
   32554: out<=0;
   32555: out<=1;
   32556: out<=1;
   32557: out<=1;
   32558: out<=0;
   32559: out<=0;
   32560: out<=1;
   32561: out<=0;
   32562: out<=0;
   32563: out<=1;
   32564: out<=1;
   32565: out<=1;
   32566: out<=1;
   32567: out<=1;
   32568: out<=0;
   32569: out<=0;
   32570: out<=1;
   32571: out<=1;
   32572: out<=0;
   32573: out<=1;
   32574: out<=0;
   32575: out<=1;
   32576: out<=1;
   32577: out<=0;
   32578: out<=1;
   32579: out<=0;
   32580: out<=1;
   32581: out<=1;
   32582: out<=0;
   32583: out<=0;
   32584: out<=1;
   32585: out<=1;
   32586: out<=1;
   32587: out<=1;
   32588: out<=1;
   32589: out<=0;
   32590: out<=0;
   32591: out<=1;
   32592: out<=1;
   32593: out<=1;
   32594: out<=0;
   32595: out<=0;
   32596: out<=0;
   32597: out<=1;
   32598: out<=0;
   32599: out<=1;
   32600: out<=0;
   32601: out<=1;
   32602: out<=1;
   32603: out<=0;
   32604: out<=1;
   32605: out<=1;
   32606: out<=1;
   32607: out<=1;
   32608: out<=1;
   32609: out<=1;
   32610: out<=1;
   32611: out<=1;
   32612: out<=0;
   32613: out<=1;
   32614: out<=1;
   32615: out<=0;
   32616: out<=1;
   32617: out<=0;
   32618: out<=1;
   32619: out<=0;
   32620: out<=0;
   32621: out<=0;
   32622: out<=1;
   32623: out<=1;
   32624: out<=1;
   32625: out<=0;
   32626: out<=0;
   32627: out<=1;
   32628: out<=1;
   32629: out<=1;
   32630: out<=1;
   32631: out<=1;
   32632: out<=0;
   32633: out<=0;
   32634: out<=1;
   32635: out<=1;
   32636: out<=0;
   32637: out<=1;
   32638: out<=0;
   32639: out<=1;
   32640: out<=0;
   32641: out<=1;
   32642: out<=0;
   32643: out<=1;
   32644: out<=0;
   32645: out<=0;
   32646: out<=1;
   32647: out<=1;
   32648: out<=0;
   32649: out<=0;
   32650: out<=0;
   32651: out<=0;
   32652: out<=0;
   32653: out<=1;
   32654: out<=1;
   32655: out<=0;
   32656: out<=0;
   32657: out<=0;
   32658: out<=1;
   32659: out<=1;
   32660: out<=1;
   32661: out<=0;
   32662: out<=1;
   32663: out<=0;
   32664: out<=1;
   32665: out<=0;
   32666: out<=0;
   32667: out<=1;
   32668: out<=0;
   32669: out<=0;
   32670: out<=0;
   32671: out<=0;
   32672: out<=1;
   32673: out<=1;
   32674: out<=1;
   32675: out<=1;
   32676: out<=0;
   32677: out<=1;
   32678: out<=1;
   32679: out<=0;
   32680: out<=1;
   32681: out<=0;
   32682: out<=1;
   32683: out<=0;
   32684: out<=0;
   32685: out<=0;
   32686: out<=1;
   32687: out<=1;
   32688: out<=1;
   32689: out<=0;
   32690: out<=0;
   32691: out<=1;
   32692: out<=1;
   32693: out<=1;
   32694: out<=1;
   32695: out<=1;
   32696: out<=0;
   32697: out<=0;
   32698: out<=1;
   32699: out<=1;
   32700: out<=0;
   32701: out<=1;
   32702: out<=0;
   32703: out<=1;
   32704: out<=0;
   32705: out<=1;
   32706: out<=0;
   32707: out<=1;
   32708: out<=0;
   32709: out<=0;
   32710: out<=1;
   32711: out<=1;
   32712: out<=0;
   32713: out<=0;
   32714: out<=0;
   32715: out<=0;
   32716: out<=0;
   32717: out<=1;
   32718: out<=1;
   32719: out<=0;
   32720: out<=1;
   32721: out<=1;
   32722: out<=0;
   32723: out<=0;
   32724: out<=0;
   32725: out<=1;
   32726: out<=0;
   32727: out<=1;
   32728: out<=0;
   32729: out<=1;
   32730: out<=1;
   32731: out<=0;
   32732: out<=1;
   32733: out<=1;
   32734: out<=1;
   32735: out<=1;
   32736: out<=0;
   32737: out<=0;
   32738: out<=0;
   32739: out<=0;
   32740: out<=1;
   32741: out<=0;
   32742: out<=0;
   32743: out<=1;
   32744: out<=0;
   32745: out<=1;
   32746: out<=0;
   32747: out<=1;
   32748: out<=1;
   32749: out<=1;
   32750: out<=0;
   32751: out<=0;
   32752: out<=1;
   32753: out<=0;
   32754: out<=0;
   32755: out<=1;
   32756: out<=1;
   32757: out<=1;
   32758: out<=1;
   32759: out<=1;
   32760: out<=0;
   32761: out<=0;
   32762: out<=1;
   32763: out<=1;
   32764: out<=0;
   32765: out<=1;
   32766: out<=0;
   32767: out<=1;
   32768: out<=0;
   32769: out<=1;
   32770: out<=0;
   32771: out<=1;
   32772: out<=0;
   32773: out<=0;
   32774: out<=1;
   32775: out<=1;
   32776: out<=0;
   32777: out<=0;
   32778: out<=0;
   32779: out<=0;
   32780: out<=0;
   32781: out<=1;
   32782: out<=1;
   32783: out<=0;
   32784: out<=1;
   32785: out<=1;
   32786: out<=0;
   32787: out<=0;
   32788: out<=0;
   32789: out<=1;
   32790: out<=0;
   32791: out<=1;
   32792: out<=0;
   32793: out<=1;
   32794: out<=1;
   32795: out<=0;
   32796: out<=1;
   32797: out<=1;
   32798: out<=1;
   32799: out<=1;
   32800: out<=0;
   32801: out<=0;
   32802: out<=0;
   32803: out<=0;
   32804: out<=1;
   32805: out<=0;
   32806: out<=0;
   32807: out<=1;
   32808: out<=0;
   32809: out<=1;
   32810: out<=0;
   32811: out<=1;
   32812: out<=1;
   32813: out<=1;
   32814: out<=0;
   32815: out<=0;
   32816: out<=1;
   32817: out<=0;
   32818: out<=0;
   32819: out<=1;
   32820: out<=1;
   32821: out<=1;
   32822: out<=1;
   32823: out<=1;
   32824: out<=0;
   32825: out<=0;
   32826: out<=1;
   32827: out<=1;
   32828: out<=0;
   32829: out<=1;
   32830: out<=0;
   32831: out<=1;
   32832: out<=0;
   32833: out<=1;
   32834: out<=0;
   32835: out<=1;
   32836: out<=0;
   32837: out<=0;
   32838: out<=1;
   32839: out<=1;
   32840: out<=0;
   32841: out<=0;
   32842: out<=0;
   32843: out<=0;
   32844: out<=0;
   32845: out<=1;
   32846: out<=1;
   32847: out<=0;
   32848: out<=0;
   32849: out<=0;
   32850: out<=1;
   32851: out<=1;
   32852: out<=1;
   32853: out<=0;
   32854: out<=1;
   32855: out<=0;
   32856: out<=1;
   32857: out<=0;
   32858: out<=0;
   32859: out<=1;
   32860: out<=0;
   32861: out<=0;
   32862: out<=0;
   32863: out<=0;
   32864: out<=1;
   32865: out<=1;
   32866: out<=1;
   32867: out<=1;
   32868: out<=0;
   32869: out<=1;
   32870: out<=1;
   32871: out<=0;
   32872: out<=1;
   32873: out<=0;
   32874: out<=1;
   32875: out<=0;
   32876: out<=0;
   32877: out<=0;
   32878: out<=1;
   32879: out<=1;
   32880: out<=1;
   32881: out<=0;
   32882: out<=0;
   32883: out<=1;
   32884: out<=1;
   32885: out<=1;
   32886: out<=1;
   32887: out<=1;
   32888: out<=0;
   32889: out<=0;
   32890: out<=1;
   32891: out<=1;
   32892: out<=0;
   32893: out<=1;
   32894: out<=0;
   32895: out<=1;
   32896: out<=0;
   32897: out<=1;
   32898: out<=0;
   32899: out<=1;
   32900: out<=0;
   32901: out<=0;
   32902: out<=1;
   32903: out<=1;
   32904: out<=0;
   32905: out<=0;
   32906: out<=0;
   32907: out<=0;
   32908: out<=0;
   32909: out<=1;
   32910: out<=1;
   32911: out<=0;
   32912: out<=0;
   32913: out<=0;
   32914: out<=1;
   32915: out<=1;
   32916: out<=1;
   32917: out<=0;
   32918: out<=1;
   32919: out<=0;
   32920: out<=1;
   32921: out<=0;
   32922: out<=0;
   32923: out<=1;
   32924: out<=0;
   32925: out<=0;
   32926: out<=0;
   32927: out<=0;
   32928: out<=0;
   32929: out<=0;
   32930: out<=0;
   32931: out<=0;
   32932: out<=1;
   32933: out<=0;
   32934: out<=0;
   32935: out<=1;
   32936: out<=0;
   32937: out<=1;
   32938: out<=0;
   32939: out<=1;
   32940: out<=1;
   32941: out<=1;
   32942: out<=0;
   32943: out<=0;
   32944: out<=0;
   32945: out<=1;
   32946: out<=1;
   32947: out<=0;
   32948: out<=0;
   32949: out<=0;
   32950: out<=0;
   32951: out<=0;
   32952: out<=1;
   32953: out<=1;
   32954: out<=0;
   32955: out<=0;
   32956: out<=1;
   32957: out<=0;
   32958: out<=1;
   32959: out<=0;
   32960: out<=0;
   32961: out<=1;
   32962: out<=0;
   32963: out<=1;
   32964: out<=0;
   32965: out<=0;
   32966: out<=1;
   32967: out<=1;
   32968: out<=0;
   32969: out<=0;
   32970: out<=0;
   32971: out<=0;
   32972: out<=0;
   32973: out<=1;
   32974: out<=1;
   32975: out<=0;
   32976: out<=1;
   32977: out<=1;
   32978: out<=0;
   32979: out<=0;
   32980: out<=0;
   32981: out<=1;
   32982: out<=0;
   32983: out<=1;
   32984: out<=0;
   32985: out<=1;
   32986: out<=1;
   32987: out<=0;
   32988: out<=1;
   32989: out<=1;
   32990: out<=1;
   32991: out<=1;
   32992: out<=1;
   32993: out<=1;
   32994: out<=1;
   32995: out<=1;
   32996: out<=0;
   32997: out<=1;
   32998: out<=1;
   32999: out<=0;
   33000: out<=1;
   33001: out<=0;
   33002: out<=1;
   33003: out<=0;
   33004: out<=0;
   33005: out<=0;
   33006: out<=1;
   33007: out<=1;
   33008: out<=0;
   33009: out<=1;
   33010: out<=1;
   33011: out<=0;
   33012: out<=0;
   33013: out<=0;
   33014: out<=0;
   33015: out<=0;
   33016: out<=1;
   33017: out<=1;
   33018: out<=0;
   33019: out<=0;
   33020: out<=1;
   33021: out<=0;
   33022: out<=1;
   33023: out<=0;
   33024: out<=0;
   33025: out<=0;
   33026: out<=1;
   33027: out<=1;
   33028: out<=1;
   33029: out<=0;
   33030: out<=1;
   33031: out<=0;
   33032: out<=1;
   33033: out<=0;
   33034: out<=0;
   33035: out<=1;
   33036: out<=0;
   33037: out<=0;
   33038: out<=0;
   33039: out<=0;
   33040: out<=0;
   33041: out<=1;
   33042: out<=0;
   33043: out<=1;
   33044: out<=0;
   33045: out<=0;
   33046: out<=1;
   33047: out<=1;
   33048: out<=0;
   33049: out<=0;
   33050: out<=0;
   33051: out<=0;
   33052: out<=0;
   33053: out<=1;
   33054: out<=1;
   33055: out<=0;
   33056: out<=1;
   33057: out<=0;
   33058: out<=0;
   33059: out<=1;
   33060: out<=1;
   33061: out<=1;
   33062: out<=1;
   33063: out<=1;
   33064: out<=0;
   33065: out<=0;
   33066: out<=1;
   33067: out<=1;
   33068: out<=0;
   33069: out<=1;
   33070: out<=0;
   33071: out<=1;
   33072: out<=1;
   33073: out<=1;
   33074: out<=1;
   33075: out<=1;
   33076: out<=0;
   33077: out<=1;
   33078: out<=1;
   33079: out<=0;
   33080: out<=1;
   33081: out<=0;
   33082: out<=1;
   33083: out<=0;
   33084: out<=0;
   33085: out<=0;
   33086: out<=1;
   33087: out<=1;
   33088: out<=1;
   33089: out<=1;
   33090: out<=0;
   33091: out<=0;
   33092: out<=0;
   33093: out<=1;
   33094: out<=0;
   33095: out<=1;
   33096: out<=0;
   33097: out<=1;
   33098: out<=1;
   33099: out<=0;
   33100: out<=1;
   33101: out<=1;
   33102: out<=1;
   33103: out<=1;
   33104: out<=0;
   33105: out<=1;
   33106: out<=0;
   33107: out<=1;
   33108: out<=0;
   33109: out<=0;
   33110: out<=1;
   33111: out<=1;
   33112: out<=0;
   33113: out<=0;
   33114: out<=0;
   33115: out<=0;
   33116: out<=0;
   33117: out<=1;
   33118: out<=1;
   33119: out<=0;
   33120: out<=1;
   33121: out<=0;
   33122: out<=0;
   33123: out<=1;
   33124: out<=1;
   33125: out<=1;
   33126: out<=1;
   33127: out<=1;
   33128: out<=0;
   33129: out<=0;
   33130: out<=1;
   33131: out<=1;
   33132: out<=0;
   33133: out<=1;
   33134: out<=0;
   33135: out<=1;
   33136: out<=0;
   33137: out<=0;
   33138: out<=0;
   33139: out<=0;
   33140: out<=1;
   33141: out<=0;
   33142: out<=0;
   33143: out<=1;
   33144: out<=0;
   33145: out<=1;
   33146: out<=0;
   33147: out<=1;
   33148: out<=1;
   33149: out<=1;
   33150: out<=0;
   33151: out<=0;
   33152: out<=1;
   33153: out<=1;
   33154: out<=0;
   33155: out<=0;
   33156: out<=0;
   33157: out<=1;
   33158: out<=0;
   33159: out<=1;
   33160: out<=0;
   33161: out<=1;
   33162: out<=1;
   33163: out<=0;
   33164: out<=1;
   33165: out<=1;
   33166: out<=1;
   33167: out<=1;
   33168: out<=0;
   33169: out<=1;
   33170: out<=0;
   33171: out<=1;
   33172: out<=0;
   33173: out<=0;
   33174: out<=1;
   33175: out<=1;
   33176: out<=0;
   33177: out<=0;
   33178: out<=0;
   33179: out<=0;
   33180: out<=0;
   33181: out<=1;
   33182: out<=1;
   33183: out<=0;
   33184: out<=0;
   33185: out<=1;
   33186: out<=1;
   33187: out<=0;
   33188: out<=0;
   33189: out<=0;
   33190: out<=0;
   33191: out<=0;
   33192: out<=1;
   33193: out<=1;
   33194: out<=0;
   33195: out<=0;
   33196: out<=1;
   33197: out<=0;
   33198: out<=1;
   33199: out<=0;
   33200: out<=1;
   33201: out<=1;
   33202: out<=1;
   33203: out<=1;
   33204: out<=0;
   33205: out<=1;
   33206: out<=1;
   33207: out<=0;
   33208: out<=1;
   33209: out<=0;
   33210: out<=1;
   33211: out<=0;
   33212: out<=0;
   33213: out<=0;
   33214: out<=1;
   33215: out<=1;
   33216: out<=0;
   33217: out<=0;
   33218: out<=1;
   33219: out<=1;
   33220: out<=1;
   33221: out<=0;
   33222: out<=1;
   33223: out<=0;
   33224: out<=1;
   33225: out<=0;
   33226: out<=0;
   33227: out<=1;
   33228: out<=0;
   33229: out<=0;
   33230: out<=0;
   33231: out<=0;
   33232: out<=0;
   33233: out<=1;
   33234: out<=0;
   33235: out<=1;
   33236: out<=0;
   33237: out<=0;
   33238: out<=1;
   33239: out<=1;
   33240: out<=0;
   33241: out<=0;
   33242: out<=0;
   33243: out<=0;
   33244: out<=0;
   33245: out<=1;
   33246: out<=1;
   33247: out<=0;
   33248: out<=0;
   33249: out<=1;
   33250: out<=1;
   33251: out<=0;
   33252: out<=0;
   33253: out<=0;
   33254: out<=0;
   33255: out<=0;
   33256: out<=1;
   33257: out<=1;
   33258: out<=0;
   33259: out<=0;
   33260: out<=1;
   33261: out<=0;
   33262: out<=1;
   33263: out<=0;
   33264: out<=0;
   33265: out<=0;
   33266: out<=0;
   33267: out<=0;
   33268: out<=1;
   33269: out<=0;
   33270: out<=0;
   33271: out<=1;
   33272: out<=0;
   33273: out<=1;
   33274: out<=0;
   33275: out<=1;
   33276: out<=1;
   33277: out<=1;
   33278: out<=0;
   33279: out<=0;
   33280: out<=0;
   33281: out<=0;
   33282: out<=0;
   33283: out<=0;
   33284: out<=1;
   33285: out<=0;
   33286: out<=0;
   33287: out<=1;
   33288: out<=0;
   33289: out<=1;
   33290: out<=0;
   33291: out<=1;
   33292: out<=1;
   33293: out<=1;
   33294: out<=0;
   33295: out<=0;
   33296: out<=0;
   33297: out<=1;
   33298: out<=1;
   33299: out<=0;
   33300: out<=0;
   33301: out<=0;
   33302: out<=0;
   33303: out<=0;
   33304: out<=1;
   33305: out<=1;
   33306: out<=0;
   33307: out<=0;
   33308: out<=1;
   33309: out<=0;
   33310: out<=1;
   33311: out<=0;
   33312: out<=0;
   33313: out<=1;
   33314: out<=0;
   33315: out<=1;
   33316: out<=0;
   33317: out<=0;
   33318: out<=1;
   33319: out<=1;
   33320: out<=0;
   33321: out<=0;
   33322: out<=0;
   33323: out<=0;
   33324: out<=0;
   33325: out<=1;
   33326: out<=1;
   33327: out<=0;
   33328: out<=0;
   33329: out<=0;
   33330: out<=1;
   33331: out<=1;
   33332: out<=1;
   33333: out<=0;
   33334: out<=1;
   33335: out<=0;
   33336: out<=1;
   33337: out<=0;
   33338: out<=0;
   33339: out<=1;
   33340: out<=0;
   33341: out<=0;
   33342: out<=0;
   33343: out<=0;
   33344: out<=1;
   33345: out<=1;
   33346: out<=1;
   33347: out<=1;
   33348: out<=0;
   33349: out<=1;
   33350: out<=1;
   33351: out<=0;
   33352: out<=1;
   33353: out<=0;
   33354: out<=1;
   33355: out<=0;
   33356: out<=0;
   33357: out<=0;
   33358: out<=1;
   33359: out<=1;
   33360: out<=0;
   33361: out<=1;
   33362: out<=1;
   33363: out<=0;
   33364: out<=0;
   33365: out<=0;
   33366: out<=0;
   33367: out<=0;
   33368: out<=1;
   33369: out<=1;
   33370: out<=0;
   33371: out<=0;
   33372: out<=1;
   33373: out<=0;
   33374: out<=1;
   33375: out<=0;
   33376: out<=0;
   33377: out<=1;
   33378: out<=0;
   33379: out<=1;
   33380: out<=0;
   33381: out<=0;
   33382: out<=1;
   33383: out<=1;
   33384: out<=0;
   33385: out<=0;
   33386: out<=0;
   33387: out<=0;
   33388: out<=0;
   33389: out<=1;
   33390: out<=1;
   33391: out<=0;
   33392: out<=1;
   33393: out<=1;
   33394: out<=0;
   33395: out<=0;
   33396: out<=0;
   33397: out<=1;
   33398: out<=0;
   33399: out<=1;
   33400: out<=0;
   33401: out<=1;
   33402: out<=1;
   33403: out<=0;
   33404: out<=1;
   33405: out<=1;
   33406: out<=1;
   33407: out<=1;
   33408: out<=0;
   33409: out<=0;
   33410: out<=0;
   33411: out<=0;
   33412: out<=1;
   33413: out<=0;
   33414: out<=0;
   33415: out<=1;
   33416: out<=0;
   33417: out<=1;
   33418: out<=0;
   33419: out<=1;
   33420: out<=1;
   33421: out<=1;
   33422: out<=0;
   33423: out<=0;
   33424: out<=1;
   33425: out<=0;
   33426: out<=0;
   33427: out<=1;
   33428: out<=1;
   33429: out<=1;
   33430: out<=1;
   33431: out<=1;
   33432: out<=0;
   33433: out<=0;
   33434: out<=1;
   33435: out<=1;
   33436: out<=0;
   33437: out<=1;
   33438: out<=0;
   33439: out<=1;
   33440: out<=0;
   33441: out<=1;
   33442: out<=0;
   33443: out<=1;
   33444: out<=0;
   33445: out<=0;
   33446: out<=1;
   33447: out<=1;
   33448: out<=0;
   33449: out<=0;
   33450: out<=0;
   33451: out<=0;
   33452: out<=0;
   33453: out<=1;
   33454: out<=1;
   33455: out<=0;
   33456: out<=1;
   33457: out<=1;
   33458: out<=0;
   33459: out<=0;
   33460: out<=0;
   33461: out<=1;
   33462: out<=0;
   33463: out<=1;
   33464: out<=0;
   33465: out<=1;
   33466: out<=1;
   33467: out<=0;
   33468: out<=1;
   33469: out<=1;
   33470: out<=1;
   33471: out<=1;
   33472: out<=1;
   33473: out<=1;
   33474: out<=1;
   33475: out<=1;
   33476: out<=0;
   33477: out<=1;
   33478: out<=1;
   33479: out<=0;
   33480: out<=1;
   33481: out<=0;
   33482: out<=1;
   33483: out<=0;
   33484: out<=0;
   33485: out<=0;
   33486: out<=1;
   33487: out<=1;
   33488: out<=1;
   33489: out<=0;
   33490: out<=0;
   33491: out<=1;
   33492: out<=1;
   33493: out<=1;
   33494: out<=1;
   33495: out<=1;
   33496: out<=0;
   33497: out<=0;
   33498: out<=1;
   33499: out<=1;
   33500: out<=0;
   33501: out<=1;
   33502: out<=0;
   33503: out<=1;
   33504: out<=0;
   33505: out<=1;
   33506: out<=0;
   33507: out<=1;
   33508: out<=0;
   33509: out<=0;
   33510: out<=1;
   33511: out<=1;
   33512: out<=0;
   33513: out<=0;
   33514: out<=0;
   33515: out<=0;
   33516: out<=0;
   33517: out<=1;
   33518: out<=1;
   33519: out<=0;
   33520: out<=0;
   33521: out<=0;
   33522: out<=1;
   33523: out<=1;
   33524: out<=1;
   33525: out<=0;
   33526: out<=1;
   33527: out<=0;
   33528: out<=1;
   33529: out<=0;
   33530: out<=0;
   33531: out<=1;
   33532: out<=0;
   33533: out<=0;
   33534: out<=0;
   33535: out<=0;
   33536: out<=0;
   33537: out<=1;
   33538: out<=1;
   33539: out<=0;
   33540: out<=0;
   33541: out<=0;
   33542: out<=0;
   33543: out<=0;
   33544: out<=1;
   33545: out<=1;
   33546: out<=0;
   33547: out<=0;
   33548: out<=1;
   33549: out<=0;
   33550: out<=1;
   33551: out<=0;
   33552: out<=1;
   33553: out<=1;
   33554: out<=1;
   33555: out<=1;
   33556: out<=0;
   33557: out<=1;
   33558: out<=1;
   33559: out<=0;
   33560: out<=1;
   33561: out<=0;
   33562: out<=1;
   33563: out<=0;
   33564: out<=0;
   33565: out<=0;
   33566: out<=1;
   33567: out<=1;
   33568: out<=1;
   33569: out<=1;
   33570: out<=0;
   33571: out<=0;
   33572: out<=0;
   33573: out<=1;
   33574: out<=0;
   33575: out<=1;
   33576: out<=0;
   33577: out<=1;
   33578: out<=1;
   33579: out<=0;
   33580: out<=1;
   33581: out<=1;
   33582: out<=1;
   33583: out<=1;
   33584: out<=0;
   33585: out<=1;
   33586: out<=0;
   33587: out<=1;
   33588: out<=0;
   33589: out<=0;
   33590: out<=1;
   33591: out<=1;
   33592: out<=0;
   33593: out<=0;
   33594: out<=0;
   33595: out<=0;
   33596: out<=0;
   33597: out<=1;
   33598: out<=1;
   33599: out<=0;
   33600: out<=0;
   33601: out<=1;
   33602: out<=1;
   33603: out<=0;
   33604: out<=0;
   33605: out<=0;
   33606: out<=0;
   33607: out<=0;
   33608: out<=1;
   33609: out<=1;
   33610: out<=0;
   33611: out<=0;
   33612: out<=1;
   33613: out<=0;
   33614: out<=1;
   33615: out<=0;
   33616: out<=0;
   33617: out<=0;
   33618: out<=0;
   33619: out<=0;
   33620: out<=1;
   33621: out<=0;
   33622: out<=0;
   33623: out<=1;
   33624: out<=0;
   33625: out<=1;
   33626: out<=0;
   33627: out<=1;
   33628: out<=1;
   33629: out<=1;
   33630: out<=0;
   33631: out<=0;
   33632: out<=0;
   33633: out<=0;
   33634: out<=1;
   33635: out<=1;
   33636: out<=1;
   33637: out<=0;
   33638: out<=1;
   33639: out<=0;
   33640: out<=1;
   33641: out<=0;
   33642: out<=0;
   33643: out<=1;
   33644: out<=0;
   33645: out<=0;
   33646: out<=0;
   33647: out<=0;
   33648: out<=0;
   33649: out<=1;
   33650: out<=0;
   33651: out<=1;
   33652: out<=0;
   33653: out<=0;
   33654: out<=1;
   33655: out<=1;
   33656: out<=0;
   33657: out<=0;
   33658: out<=0;
   33659: out<=0;
   33660: out<=0;
   33661: out<=1;
   33662: out<=1;
   33663: out<=0;
   33664: out<=1;
   33665: out<=0;
   33666: out<=0;
   33667: out<=1;
   33668: out<=1;
   33669: out<=1;
   33670: out<=1;
   33671: out<=1;
   33672: out<=0;
   33673: out<=0;
   33674: out<=1;
   33675: out<=1;
   33676: out<=0;
   33677: out<=1;
   33678: out<=0;
   33679: out<=1;
   33680: out<=1;
   33681: out<=1;
   33682: out<=1;
   33683: out<=1;
   33684: out<=0;
   33685: out<=1;
   33686: out<=1;
   33687: out<=0;
   33688: out<=1;
   33689: out<=0;
   33690: out<=1;
   33691: out<=0;
   33692: out<=0;
   33693: out<=0;
   33694: out<=1;
   33695: out<=1;
   33696: out<=0;
   33697: out<=0;
   33698: out<=1;
   33699: out<=1;
   33700: out<=1;
   33701: out<=0;
   33702: out<=1;
   33703: out<=0;
   33704: out<=1;
   33705: out<=0;
   33706: out<=0;
   33707: out<=1;
   33708: out<=0;
   33709: out<=0;
   33710: out<=0;
   33711: out<=0;
   33712: out<=0;
   33713: out<=1;
   33714: out<=0;
   33715: out<=1;
   33716: out<=0;
   33717: out<=0;
   33718: out<=1;
   33719: out<=1;
   33720: out<=0;
   33721: out<=0;
   33722: out<=0;
   33723: out<=0;
   33724: out<=0;
   33725: out<=1;
   33726: out<=1;
   33727: out<=0;
   33728: out<=1;
   33729: out<=0;
   33730: out<=0;
   33731: out<=1;
   33732: out<=1;
   33733: out<=1;
   33734: out<=1;
   33735: out<=1;
   33736: out<=0;
   33737: out<=0;
   33738: out<=1;
   33739: out<=1;
   33740: out<=0;
   33741: out<=1;
   33742: out<=0;
   33743: out<=1;
   33744: out<=0;
   33745: out<=0;
   33746: out<=0;
   33747: out<=0;
   33748: out<=1;
   33749: out<=0;
   33750: out<=0;
   33751: out<=1;
   33752: out<=0;
   33753: out<=1;
   33754: out<=0;
   33755: out<=1;
   33756: out<=1;
   33757: out<=1;
   33758: out<=0;
   33759: out<=0;
   33760: out<=1;
   33761: out<=1;
   33762: out<=0;
   33763: out<=0;
   33764: out<=0;
   33765: out<=1;
   33766: out<=0;
   33767: out<=1;
   33768: out<=0;
   33769: out<=1;
   33770: out<=1;
   33771: out<=0;
   33772: out<=1;
   33773: out<=1;
   33774: out<=1;
   33775: out<=1;
   33776: out<=0;
   33777: out<=1;
   33778: out<=0;
   33779: out<=1;
   33780: out<=0;
   33781: out<=0;
   33782: out<=1;
   33783: out<=1;
   33784: out<=0;
   33785: out<=0;
   33786: out<=0;
   33787: out<=0;
   33788: out<=0;
   33789: out<=1;
   33790: out<=1;
   33791: out<=0;
   33792: out<=0;
   33793: out<=0;
   33794: out<=1;
   33795: out<=1;
   33796: out<=0;
   33797: out<=1;
   33798: out<=0;
   33799: out<=1;
   33800: out<=0;
   33801: out<=1;
   33802: out<=1;
   33803: out<=0;
   33804: out<=0;
   33805: out<=0;
   33806: out<=0;
   33807: out<=0;
   33808: out<=1;
   33809: out<=0;
   33810: out<=1;
   33811: out<=0;
   33812: out<=0;
   33813: out<=0;
   33814: out<=1;
   33815: out<=1;
   33816: out<=0;
   33817: out<=0;
   33818: out<=0;
   33819: out<=0;
   33820: out<=1;
   33821: out<=0;
   33822: out<=0;
   33823: out<=1;
   33824: out<=0;
   33825: out<=1;
   33826: out<=1;
   33827: out<=0;
   33828: out<=1;
   33829: out<=1;
   33830: out<=1;
   33831: out<=1;
   33832: out<=0;
   33833: out<=0;
   33834: out<=1;
   33835: out<=1;
   33836: out<=1;
   33837: out<=0;
   33838: out<=1;
   33839: out<=0;
   33840: out<=1;
   33841: out<=1;
   33842: out<=1;
   33843: out<=1;
   33844: out<=1;
   33845: out<=0;
   33846: out<=0;
   33847: out<=1;
   33848: out<=0;
   33849: out<=1;
   33850: out<=0;
   33851: out<=1;
   33852: out<=0;
   33853: out<=0;
   33854: out<=1;
   33855: out<=1;
   33856: out<=1;
   33857: out<=1;
   33858: out<=0;
   33859: out<=0;
   33860: out<=1;
   33861: out<=0;
   33862: out<=1;
   33863: out<=0;
   33864: out<=1;
   33865: out<=0;
   33866: out<=0;
   33867: out<=1;
   33868: out<=1;
   33869: out<=1;
   33870: out<=1;
   33871: out<=1;
   33872: out<=1;
   33873: out<=0;
   33874: out<=1;
   33875: out<=0;
   33876: out<=0;
   33877: out<=0;
   33878: out<=1;
   33879: out<=1;
   33880: out<=0;
   33881: out<=0;
   33882: out<=0;
   33883: out<=0;
   33884: out<=1;
   33885: out<=0;
   33886: out<=0;
   33887: out<=1;
   33888: out<=0;
   33889: out<=1;
   33890: out<=1;
   33891: out<=0;
   33892: out<=1;
   33893: out<=1;
   33894: out<=1;
   33895: out<=1;
   33896: out<=0;
   33897: out<=0;
   33898: out<=1;
   33899: out<=1;
   33900: out<=1;
   33901: out<=0;
   33902: out<=1;
   33903: out<=0;
   33904: out<=0;
   33905: out<=0;
   33906: out<=0;
   33907: out<=0;
   33908: out<=0;
   33909: out<=1;
   33910: out<=1;
   33911: out<=0;
   33912: out<=1;
   33913: out<=0;
   33914: out<=1;
   33915: out<=0;
   33916: out<=1;
   33917: out<=1;
   33918: out<=0;
   33919: out<=0;
   33920: out<=1;
   33921: out<=1;
   33922: out<=0;
   33923: out<=0;
   33924: out<=1;
   33925: out<=0;
   33926: out<=1;
   33927: out<=0;
   33928: out<=1;
   33929: out<=0;
   33930: out<=0;
   33931: out<=1;
   33932: out<=1;
   33933: out<=1;
   33934: out<=1;
   33935: out<=1;
   33936: out<=1;
   33937: out<=0;
   33938: out<=1;
   33939: out<=0;
   33940: out<=0;
   33941: out<=0;
   33942: out<=1;
   33943: out<=1;
   33944: out<=0;
   33945: out<=0;
   33946: out<=0;
   33947: out<=0;
   33948: out<=1;
   33949: out<=0;
   33950: out<=0;
   33951: out<=1;
   33952: out<=1;
   33953: out<=0;
   33954: out<=0;
   33955: out<=1;
   33956: out<=0;
   33957: out<=0;
   33958: out<=0;
   33959: out<=0;
   33960: out<=1;
   33961: out<=1;
   33962: out<=0;
   33963: out<=0;
   33964: out<=0;
   33965: out<=1;
   33966: out<=0;
   33967: out<=1;
   33968: out<=1;
   33969: out<=1;
   33970: out<=1;
   33971: out<=1;
   33972: out<=1;
   33973: out<=0;
   33974: out<=0;
   33975: out<=1;
   33976: out<=0;
   33977: out<=1;
   33978: out<=0;
   33979: out<=1;
   33980: out<=0;
   33981: out<=0;
   33982: out<=1;
   33983: out<=1;
   33984: out<=0;
   33985: out<=0;
   33986: out<=1;
   33987: out<=1;
   33988: out<=0;
   33989: out<=1;
   33990: out<=0;
   33991: out<=1;
   33992: out<=0;
   33993: out<=1;
   33994: out<=1;
   33995: out<=0;
   33996: out<=0;
   33997: out<=0;
   33998: out<=0;
   33999: out<=0;
   34000: out<=1;
   34001: out<=0;
   34002: out<=1;
   34003: out<=0;
   34004: out<=0;
   34005: out<=0;
   34006: out<=1;
   34007: out<=1;
   34008: out<=0;
   34009: out<=0;
   34010: out<=0;
   34011: out<=0;
   34012: out<=1;
   34013: out<=0;
   34014: out<=0;
   34015: out<=1;
   34016: out<=1;
   34017: out<=0;
   34018: out<=0;
   34019: out<=1;
   34020: out<=0;
   34021: out<=0;
   34022: out<=0;
   34023: out<=0;
   34024: out<=1;
   34025: out<=1;
   34026: out<=0;
   34027: out<=0;
   34028: out<=0;
   34029: out<=1;
   34030: out<=0;
   34031: out<=1;
   34032: out<=0;
   34033: out<=0;
   34034: out<=0;
   34035: out<=0;
   34036: out<=0;
   34037: out<=1;
   34038: out<=1;
   34039: out<=0;
   34040: out<=1;
   34041: out<=0;
   34042: out<=1;
   34043: out<=0;
   34044: out<=1;
   34045: out<=1;
   34046: out<=0;
   34047: out<=0;
   34048: out<=1;
   34049: out<=0;
   34050: out<=1;
   34051: out<=0;
   34052: out<=0;
   34053: out<=0;
   34054: out<=1;
   34055: out<=1;
   34056: out<=0;
   34057: out<=0;
   34058: out<=0;
   34059: out<=0;
   34060: out<=1;
   34061: out<=0;
   34062: out<=0;
   34063: out<=1;
   34064: out<=1;
   34065: out<=1;
   34066: out<=0;
   34067: out<=0;
   34068: out<=1;
   34069: out<=0;
   34070: out<=1;
   34071: out<=0;
   34072: out<=1;
   34073: out<=0;
   34074: out<=0;
   34075: out<=1;
   34076: out<=1;
   34077: out<=1;
   34078: out<=1;
   34079: out<=1;
   34080: out<=0;
   34081: out<=0;
   34082: out<=0;
   34083: out<=0;
   34084: out<=0;
   34085: out<=1;
   34086: out<=1;
   34087: out<=0;
   34088: out<=1;
   34089: out<=0;
   34090: out<=1;
   34091: out<=0;
   34092: out<=1;
   34093: out<=1;
   34094: out<=0;
   34095: out<=0;
   34096: out<=0;
   34097: out<=1;
   34098: out<=1;
   34099: out<=0;
   34100: out<=1;
   34101: out<=1;
   34102: out<=1;
   34103: out<=1;
   34104: out<=0;
   34105: out<=0;
   34106: out<=1;
   34107: out<=1;
   34108: out<=1;
   34109: out<=0;
   34110: out<=1;
   34111: out<=0;
   34112: out<=1;
   34113: out<=0;
   34114: out<=1;
   34115: out<=0;
   34116: out<=0;
   34117: out<=0;
   34118: out<=1;
   34119: out<=1;
   34120: out<=0;
   34121: out<=0;
   34122: out<=0;
   34123: out<=0;
   34124: out<=1;
   34125: out<=0;
   34126: out<=0;
   34127: out<=1;
   34128: out<=0;
   34129: out<=0;
   34130: out<=1;
   34131: out<=1;
   34132: out<=0;
   34133: out<=1;
   34134: out<=0;
   34135: out<=1;
   34136: out<=0;
   34137: out<=1;
   34138: out<=1;
   34139: out<=0;
   34140: out<=0;
   34141: out<=0;
   34142: out<=0;
   34143: out<=0;
   34144: out<=1;
   34145: out<=1;
   34146: out<=1;
   34147: out<=1;
   34148: out<=1;
   34149: out<=0;
   34150: out<=0;
   34151: out<=1;
   34152: out<=0;
   34153: out<=1;
   34154: out<=0;
   34155: out<=1;
   34156: out<=0;
   34157: out<=0;
   34158: out<=1;
   34159: out<=1;
   34160: out<=0;
   34161: out<=1;
   34162: out<=1;
   34163: out<=0;
   34164: out<=1;
   34165: out<=1;
   34166: out<=1;
   34167: out<=1;
   34168: out<=0;
   34169: out<=0;
   34170: out<=1;
   34171: out<=1;
   34172: out<=1;
   34173: out<=0;
   34174: out<=1;
   34175: out<=0;
   34176: out<=1;
   34177: out<=0;
   34178: out<=1;
   34179: out<=0;
   34180: out<=0;
   34181: out<=0;
   34182: out<=1;
   34183: out<=1;
   34184: out<=0;
   34185: out<=0;
   34186: out<=0;
   34187: out<=0;
   34188: out<=1;
   34189: out<=0;
   34190: out<=0;
   34191: out<=1;
   34192: out<=0;
   34193: out<=0;
   34194: out<=1;
   34195: out<=1;
   34196: out<=0;
   34197: out<=1;
   34198: out<=0;
   34199: out<=1;
   34200: out<=0;
   34201: out<=1;
   34202: out<=1;
   34203: out<=0;
   34204: out<=0;
   34205: out<=0;
   34206: out<=0;
   34207: out<=0;
   34208: out<=0;
   34209: out<=0;
   34210: out<=0;
   34211: out<=0;
   34212: out<=0;
   34213: out<=1;
   34214: out<=1;
   34215: out<=0;
   34216: out<=1;
   34217: out<=0;
   34218: out<=1;
   34219: out<=0;
   34220: out<=1;
   34221: out<=1;
   34222: out<=0;
   34223: out<=0;
   34224: out<=1;
   34225: out<=0;
   34226: out<=0;
   34227: out<=1;
   34228: out<=0;
   34229: out<=0;
   34230: out<=0;
   34231: out<=0;
   34232: out<=1;
   34233: out<=1;
   34234: out<=0;
   34235: out<=0;
   34236: out<=0;
   34237: out<=1;
   34238: out<=0;
   34239: out<=1;
   34240: out<=1;
   34241: out<=0;
   34242: out<=1;
   34243: out<=0;
   34244: out<=0;
   34245: out<=0;
   34246: out<=1;
   34247: out<=1;
   34248: out<=0;
   34249: out<=0;
   34250: out<=0;
   34251: out<=0;
   34252: out<=1;
   34253: out<=0;
   34254: out<=0;
   34255: out<=1;
   34256: out<=1;
   34257: out<=1;
   34258: out<=0;
   34259: out<=0;
   34260: out<=1;
   34261: out<=0;
   34262: out<=1;
   34263: out<=0;
   34264: out<=1;
   34265: out<=0;
   34266: out<=0;
   34267: out<=1;
   34268: out<=1;
   34269: out<=1;
   34270: out<=1;
   34271: out<=1;
   34272: out<=1;
   34273: out<=1;
   34274: out<=1;
   34275: out<=1;
   34276: out<=1;
   34277: out<=0;
   34278: out<=0;
   34279: out<=1;
   34280: out<=0;
   34281: out<=1;
   34282: out<=0;
   34283: out<=1;
   34284: out<=0;
   34285: out<=0;
   34286: out<=1;
   34287: out<=1;
   34288: out<=1;
   34289: out<=0;
   34290: out<=0;
   34291: out<=1;
   34292: out<=0;
   34293: out<=0;
   34294: out<=0;
   34295: out<=0;
   34296: out<=1;
   34297: out<=1;
   34298: out<=0;
   34299: out<=0;
   34300: out<=0;
   34301: out<=1;
   34302: out<=0;
   34303: out<=1;
   34304: out<=1;
   34305: out<=0;
   34306: out<=0;
   34307: out<=1;
   34308: out<=0;
   34309: out<=0;
   34310: out<=0;
   34311: out<=0;
   34312: out<=1;
   34313: out<=1;
   34314: out<=0;
   34315: out<=0;
   34316: out<=0;
   34317: out<=1;
   34318: out<=0;
   34319: out<=1;
   34320: out<=1;
   34321: out<=1;
   34322: out<=1;
   34323: out<=1;
   34324: out<=1;
   34325: out<=0;
   34326: out<=0;
   34327: out<=1;
   34328: out<=0;
   34329: out<=1;
   34330: out<=0;
   34331: out<=1;
   34332: out<=0;
   34333: out<=0;
   34334: out<=1;
   34335: out<=1;
   34336: out<=1;
   34337: out<=1;
   34338: out<=0;
   34339: out<=0;
   34340: out<=1;
   34341: out<=0;
   34342: out<=1;
   34343: out<=0;
   34344: out<=1;
   34345: out<=0;
   34346: out<=0;
   34347: out<=1;
   34348: out<=1;
   34349: out<=1;
   34350: out<=1;
   34351: out<=1;
   34352: out<=1;
   34353: out<=0;
   34354: out<=1;
   34355: out<=0;
   34356: out<=0;
   34357: out<=0;
   34358: out<=1;
   34359: out<=1;
   34360: out<=0;
   34361: out<=0;
   34362: out<=0;
   34363: out<=0;
   34364: out<=1;
   34365: out<=0;
   34366: out<=0;
   34367: out<=1;
   34368: out<=1;
   34369: out<=0;
   34370: out<=0;
   34371: out<=1;
   34372: out<=0;
   34373: out<=0;
   34374: out<=0;
   34375: out<=0;
   34376: out<=1;
   34377: out<=1;
   34378: out<=0;
   34379: out<=0;
   34380: out<=0;
   34381: out<=1;
   34382: out<=0;
   34383: out<=1;
   34384: out<=0;
   34385: out<=0;
   34386: out<=0;
   34387: out<=0;
   34388: out<=0;
   34389: out<=1;
   34390: out<=1;
   34391: out<=0;
   34392: out<=1;
   34393: out<=0;
   34394: out<=1;
   34395: out<=0;
   34396: out<=1;
   34397: out<=1;
   34398: out<=0;
   34399: out<=0;
   34400: out<=0;
   34401: out<=0;
   34402: out<=1;
   34403: out<=1;
   34404: out<=0;
   34405: out<=1;
   34406: out<=0;
   34407: out<=1;
   34408: out<=0;
   34409: out<=1;
   34410: out<=1;
   34411: out<=0;
   34412: out<=0;
   34413: out<=0;
   34414: out<=0;
   34415: out<=0;
   34416: out<=1;
   34417: out<=0;
   34418: out<=1;
   34419: out<=0;
   34420: out<=0;
   34421: out<=0;
   34422: out<=1;
   34423: out<=1;
   34424: out<=0;
   34425: out<=0;
   34426: out<=0;
   34427: out<=0;
   34428: out<=1;
   34429: out<=0;
   34430: out<=0;
   34431: out<=1;
   34432: out<=0;
   34433: out<=1;
   34434: out<=1;
   34435: out<=0;
   34436: out<=1;
   34437: out<=1;
   34438: out<=1;
   34439: out<=1;
   34440: out<=0;
   34441: out<=0;
   34442: out<=1;
   34443: out<=1;
   34444: out<=1;
   34445: out<=0;
   34446: out<=1;
   34447: out<=0;
   34448: out<=1;
   34449: out<=1;
   34450: out<=1;
   34451: out<=1;
   34452: out<=1;
   34453: out<=0;
   34454: out<=0;
   34455: out<=1;
   34456: out<=0;
   34457: out<=1;
   34458: out<=0;
   34459: out<=1;
   34460: out<=0;
   34461: out<=0;
   34462: out<=1;
   34463: out<=1;
   34464: out<=0;
   34465: out<=0;
   34466: out<=1;
   34467: out<=1;
   34468: out<=0;
   34469: out<=1;
   34470: out<=0;
   34471: out<=1;
   34472: out<=0;
   34473: out<=1;
   34474: out<=1;
   34475: out<=0;
   34476: out<=0;
   34477: out<=0;
   34478: out<=0;
   34479: out<=0;
   34480: out<=1;
   34481: out<=0;
   34482: out<=1;
   34483: out<=0;
   34484: out<=0;
   34485: out<=0;
   34486: out<=1;
   34487: out<=1;
   34488: out<=0;
   34489: out<=0;
   34490: out<=0;
   34491: out<=0;
   34492: out<=1;
   34493: out<=0;
   34494: out<=0;
   34495: out<=1;
   34496: out<=0;
   34497: out<=1;
   34498: out<=1;
   34499: out<=0;
   34500: out<=1;
   34501: out<=1;
   34502: out<=1;
   34503: out<=1;
   34504: out<=0;
   34505: out<=0;
   34506: out<=1;
   34507: out<=1;
   34508: out<=1;
   34509: out<=0;
   34510: out<=1;
   34511: out<=0;
   34512: out<=0;
   34513: out<=0;
   34514: out<=0;
   34515: out<=0;
   34516: out<=0;
   34517: out<=1;
   34518: out<=1;
   34519: out<=0;
   34520: out<=1;
   34521: out<=0;
   34522: out<=1;
   34523: out<=0;
   34524: out<=1;
   34525: out<=1;
   34526: out<=0;
   34527: out<=0;
   34528: out<=1;
   34529: out<=1;
   34530: out<=0;
   34531: out<=0;
   34532: out<=1;
   34533: out<=0;
   34534: out<=1;
   34535: out<=0;
   34536: out<=1;
   34537: out<=0;
   34538: out<=0;
   34539: out<=1;
   34540: out<=1;
   34541: out<=1;
   34542: out<=1;
   34543: out<=1;
   34544: out<=1;
   34545: out<=0;
   34546: out<=1;
   34547: out<=0;
   34548: out<=0;
   34549: out<=0;
   34550: out<=1;
   34551: out<=1;
   34552: out<=0;
   34553: out<=0;
   34554: out<=0;
   34555: out<=0;
   34556: out<=1;
   34557: out<=0;
   34558: out<=0;
   34559: out<=1;
   34560: out<=0;
   34561: out<=0;
   34562: out<=0;
   34563: out<=0;
   34564: out<=0;
   34565: out<=1;
   34566: out<=1;
   34567: out<=0;
   34568: out<=1;
   34569: out<=0;
   34570: out<=1;
   34571: out<=0;
   34572: out<=1;
   34573: out<=1;
   34574: out<=0;
   34575: out<=0;
   34576: out<=1;
   34577: out<=0;
   34578: out<=0;
   34579: out<=1;
   34580: out<=0;
   34581: out<=0;
   34582: out<=0;
   34583: out<=0;
   34584: out<=1;
   34585: out<=1;
   34586: out<=0;
   34587: out<=0;
   34588: out<=0;
   34589: out<=1;
   34590: out<=0;
   34591: out<=1;
   34592: out<=1;
   34593: out<=0;
   34594: out<=1;
   34595: out<=0;
   34596: out<=0;
   34597: out<=0;
   34598: out<=1;
   34599: out<=1;
   34600: out<=0;
   34601: out<=0;
   34602: out<=0;
   34603: out<=0;
   34604: out<=1;
   34605: out<=0;
   34606: out<=0;
   34607: out<=1;
   34608: out<=0;
   34609: out<=0;
   34610: out<=1;
   34611: out<=1;
   34612: out<=0;
   34613: out<=1;
   34614: out<=0;
   34615: out<=1;
   34616: out<=0;
   34617: out<=1;
   34618: out<=1;
   34619: out<=0;
   34620: out<=0;
   34621: out<=0;
   34622: out<=0;
   34623: out<=0;
   34624: out<=1;
   34625: out<=1;
   34626: out<=1;
   34627: out<=1;
   34628: out<=1;
   34629: out<=0;
   34630: out<=0;
   34631: out<=1;
   34632: out<=0;
   34633: out<=1;
   34634: out<=0;
   34635: out<=1;
   34636: out<=0;
   34637: out<=0;
   34638: out<=1;
   34639: out<=1;
   34640: out<=1;
   34641: out<=0;
   34642: out<=0;
   34643: out<=1;
   34644: out<=0;
   34645: out<=0;
   34646: out<=0;
   34647: out<=0;
   34648: out<=1;
   34649: out<=1;
   34650: out<=0;
   34651: out<=0;
   34652: out<=0;
   34653: out<=1;
   34654: out<=0;
   34655: out<=1;
   34656: out<=1;
   34657: out<=0;
   34658: out<=1;
   34659: out<=0;
   34660: out<=0;
   34661: out<=0;
   34662: out<=1;
   34663: out<=1;
   34664: out<=0;
   34665: out<=0;
   34666: out<=0;
   34667: out<=0;
   34668: out<=1;
   34669: out<=0;
   34670: out<=0;
   34671: out<=1;
   34672: out<=1;
   34673: out<=1;
   34674: out<=0;
   34675: out<=0;
   34676: out<=1;
   34677: out<=0;
   34678: out<=1;
   34679: out<=0;
   34680: out<=1;
   34681: out<=0;
   34682: out<=0;
   34683: out<=1;
   34684: out<=1;
   34685: out<=1;
   34686: out<=1;
   34687: out<=1;
   34688: out<=0;
   34689: out<=0;
   34690: out<=0;
   34691: out<=0;
   34692: out<=0;
   34693: out<=1;
   34694: out<=1;
   34695: out<=0;
   34696: out<=1;
   34697: out<=0;
   34698: out<=1;
   34699: out<=0;
   34700: out<=1;
   34701: out<=1;
   34702: out<=0;
   34703: out<=0;
   34704: out<=0;
   34705: out<=1;
   34706: out<=1;
   34707: out<=0;
   34708: out<=1;
   34709: out<=1;
   34710: out<=1;
   34711: out<=1;
   34712: out<=0;
   34713: out<=0;
   34714: out<=1;
   34715: out<=1;
   34716: out<=1;
   34717: out<=0;
   34718: out<=1;
   34719: out<=0;
   34720: out<=1;
   34721: out<=0;
   34722: out<=1;
   34723: out<=0;
   34724: out<=0;
   34725: out<=0;
   34726: out<=1;
   34727: out<=1;
   34728: out<=0;
   34729: out<=0;
   34730: out<=0;
   34731: out<=0;
   34732: out<=1;
   34733: out<=0;
   34734: out<=0;
   34735: out<=1;
   34736: out<=1;
   34737: out<=1;
   34738: out<=0;
   34739: out<=0;
   34740: out<=1;
   34741: out<=0;
   34742: out<=1;
   34743: out<=0;
   34744: out<=1;
   34745: out<=0;
   34746: out<=0;
   34747: out<=1;
   34748: out<=1;
   34749: out<=1;
   34750: out<=1;
   34751: out<=1;
   34752: out<=1;
   34753: out<=1;
   34754: out<=1;
   34755: out<=1;
   34756: out<=1;
   34757: out<=0;
   34758: out<=0;
   34759: out<=1;
   34760: out<=0;
   34761: out<=1;
   34762: out<=0;
   34763: out<=1;
   34764: out<=0;
   34765: out<=0;
   34766: out<=1;
   34767: out<=1;
   34768: out<=0;
   34769: out<=1;
   34770: out<=1;
   34771: out<=0;
   34772: out<=1;
   34773: out<=1;
   34774: out<=1;
   34775: out<=1;
   34776: out<=0;
   34777: out<=0;
   34778: out<=1;
   34779: out<=1;
   34780: out<=1;
   34781: out<=0;
   34782: out<=1;
   34783: out<=0;
   34784: out<=1;
   34785: out<=0;
   34786: out<=1;
   34787: out<=0;
   34788: out<=0;
   34789: out<=0;
   34790: out<=1;
   34791: out<=1;
   34792: out<=0;
   34793: out<=0;
   34794: out<=0;
   34795: out<=0;
   34796: out<=1;
   34797: out<=0;
   34798: out<=0;
   34799: out<=1;
   34800: out<=0;
   34801: out<=0;
   34802: out<=1;
   34803: out<=1;
   34804: out<=0;
   34805: out<=1;
   34806: out<=0;
   34807: out<=1;
   34808: out<=0;
   34809: out<=1;
   34810: out<=1;
   34811: out<=0;
   34812: out<=0;
   34813: out<=0;
   34814: out<=0;
   34815: out<=0;
   34816: out<=0;
   34817: out<=0;
   34818: out<=0;
   34819: out<=0;
   34820: out<=0;
   34821: out<=1;
   34822: out<=1;
   34823: out<=0;
   34824: out<=0;
   34825: out<=1;
   34826: out<=0;
   34827: out<=1;
   34828: out<=0;
   34829: out<=0;
   34830: out<=1;
   34831: out<=1;
   34832: out<=1;
   34833: out<=0;
   34834: out<=0;
   34835: out<=1;
   34836: out<=0;
   34837: out<=0;
   34838: out<=0;
   34839: out<=0;
   34840: out<=0;
   34841: out<=0;
   34842: out<=1;
   34843: out<=1;
   34844: out<=1;
   34845: out<=0;
   34846: out<=1;
   34847: out<=0;
   34848: out<=0;
   34849: out<=1;
   34850: out<=0;
   34851: out<=1;
   34852: out<=1;
   34853: out<=1;
   34854: out<=0;
   34855: out<=0;
   34856: out<=0;
   34857: out<=0;
   34858: out<=0;
   34859: out<=0;
   34860: out<=1;
   34861: out<=0;
   34862: out<=0;
   34863: out<=1;
   34864: out<=1;
   34865: out<=1;
   34866: out<=0;
   34867: out<=0;
   34868: out<=1;
   34869: out<=0;
   34870: out<=1;
   34871: out<=0;
   34872: out<=0;
   34873: out<=1;
   34874: out<=1;
   34875: out<=0;
   34876: out<=0;
   34877: out<=0;
   34878: out<=0;
   34879: out<=0;
   34880: out<=1;
   34881: out<=1;
   34882: out<=1;
   34883: out<=1;
   34884: out<=1;
   34885: out<=0;
   34886: out<=0;
   34887: out<=1;
   34888: out<=1;
   34889: out<=0;
   34890: out<=1;
   34891: out<=0;
   34892: out<=1;
   34893: out<=1;
   34894: out<=0;
   34895: out<=0;
   34896: out<=1;
   34897: out<=0;
   34898: out<=0;
   34899: out<=1;
   34900: out<=0;
   34901: out<=0;
   34902: out<=0;
   34903: out<=0;
   34904: out<=0;
   34905: out<=0;
   34906: out<=1;
   34907: out<=1;
   34908: out<=1;
   34909: out<=0;
   34910: out<=1;
   34911: out<=0;
   34912: out<=0;
   34913: out<=1;
   34914: out<=0;
   34915: out<=1;
   34916: out<=1;
   34917: out<=1;
   34918: out<=0;
   34919: out<=0;
   34920: out<=0;
   34921: out<=0;
   34922: out<=0;
   34923: out<=0;
   34924: out<=1;
   34925: out<=0;
   34926: out<=0;
   34927: out<=1;
   34928: out<=0;
   34929: out<=0;
   34930: out<=1;
   34931: out<=1;
   34932: out<=0;
   34933: out<=1;
   34934: out<=0;
   34935: out<=1;
   34936: out<=1;
   34937: out<=0;
   34938: out<=0;
   34939: out<=1;
   34940: out<=1;
   34941: out<=1;
   34942: out<=1;
   34943: out<=1;
   34944: out<=0;
   34945: out<=0;
   34946: out<=0;
   34947: out<=0;
   34948: out<=0;
   34949: out<=1;
   34950: out<=1;
   34951: out<=0;
   34952: out<=0;
   34953: out<=1;
   34954: out<=0;
   34955: out<=1;
   34956: out<=0;
   34957: out<=0;
   34958: out<=1;
   34959: out<=1;
   34960: out<=0;
   34961: out<=1;
   34962: out<=1;
   34963: out<=0;
   34964: out<=1;
   34965: out<=1;
   34966: out<=1;
   34967: out<=1;
   34968: out<=1;
   34969: out<=1;
   34970: out<=0;
   34971: out<=0;
   34972: out<=0;
   34973: out<=1;
   34974: out<=0;
   34975: out<=1;
   34976: out<=0;
   34977: out<=1;
   34978: out<=0;
   34979: out<=1;
   34980: out<=1;
   34981: out<=1;
   34982: out<=0;
   34983: out<=0;
   34984: out<=0;
   34985: out<=0;
   34986: out<=0;
   34987: out<=0;
   34988: out<=1;
   34989: out<=0;
   34990: out<=0;
   34991: out<=1;
   34992: out<=0;
   34993: out<=0;
   34994: out<=1;
   34995: out<=1;
   34996: out<=0;
   34997: out<=1;
   34998: out<=0;
   34999: out<=1;
   35000: out<=1;
   35001: out<=0;
   35002: out<=0;
   35003: out<=1;
   35004: out<=1;
   35005: out<=1;
   35006: out<=1;
   35007: out<=1;
   35008: out<=1;
   35009: out<=1;
   35010: out<=1;
   35011: out<=1;
   35012: out<=1;
   35013: out<=0;
   35014: out<=0;
   35015: out<=1;
   35016: out<=1;
   35017: out<=0;
   35018: out<=1;
   35019: out<=0;
   35020: out<=1;
   35021: out<=1;
   35022: out<=0;
   35023: out<=0;
   35024: out<=0;
   35025: out<=1;
   35026: out<=1;
   35027: out<=0;
   35028: out<=1;
   35029: out<=1;
   35030: out<=1;
   35031: out<=1;
   35032: out<=1;
   35033: out<=1;
   35034: out<=0;
   35035: out<=0;
   35036: out<=0;
   35037: out<=1;
   35038: out<=0;
   35039: out<=1;
   35040: out<=0;
   35041: out<=1;
   35042: out<=0;
   35043: out<=1;
   35044: out<=1;
   35045: out<=1;
   35046: out<=0;
   35047: out<=0;
   35048: out<=0;
   35049: out<=0;
   35050: out<=0;
   35051: out<=0;
   35052: out<=1;
   35053: out<=0;
   35054: out<=0;
   35055: out<=1;
   35056: out<=1;
   35057: out<=1;
   35058: out<=0;
   35059: out<=0;
   35060: out<=1;
   35061: out<=0;
   35062: out<=1;
   35063: out<=0;
   35064: out<=0;
   35065: out<=1;
   35066: out<=1;
   35067: out<=0;
   35068: out<=0;
   35069: out<=0;
   35070: out<=0;
   35071: out<=0;
   35072: out<=1;
   35073: out<=0;
   35074: out<=0;
   35075: out<=1;
   35076: out<=0;
   35077: out<=0;
   35078: out<=0;
   35079: out<=0;
   35080: out<=0;
   35081: out<=0;
   35082: out<=1;
   35083: out<=1;
   35084: out<=1;
   35085: out<=0;
   35086: out<=1;
   35087: out<=0;
   35088: out<=1;
   35089: out<=1;
   35090: out<=1;
   35091: out<=1;
   35092: out<=1;
   35093: out<=0;
   35094: out<=0;
   35095: out<=1;
   35096: out<=1;
   35097: out<=0;
   35098: out<=1;
   35099: out<=0;
   35100: out<=1;
   35101: out<=1;
   35102: out<=0;
   35103: out<=0;
   35104: out<=0;
   35105: out<=0;
   35106: out<=1;
   35107: out<=1;
   35108: out<=0;
   35109: out<=1;
   35110: out<=0;
   35111: out<=1;
   35112: out<=1;
   35113: out<=0;
   35114: out<=0;
   35115: out<=1;
   35116: out<=1;
   35117: out<=1;
   35118: out<=1;
   35119: out<=1;
   35120: out<=0;
   35121: out<=1;
   35122: out<=0;
   35123: out<=1;
   35124: out<=1;
   35125: out<=1;
   35126: out<=0;
   35127: out<=0;
   35128: out<=0;
   35129: out<=0;
   35130: out<=0;
   35131: out<=0;
   35132: out<=1;
   35133: out<=0;
   35134: out<=0;
   35135: out<=1;
   35136: out<=1;
   35137: out<=0;
   35138: out<=0;
   35139: out<=1;
   35140: out<=0;
   35141: out<=0;
   35142: out<=0;
   35143: out<=0;
   35144: out<=0;
   35145: out<=0;
   35146: out<=1;
   35147: out<=1;
   35148: out<=1;
   35149: out<=0;
   35150: out<=1;
   35151: out<=0;
   35152: out<=0;
   35153: out<=0;
   35154: out<=0;
   35155: out<=0;
   35156: out<=0;
   35157: out<=1;
   35158: out<=1;
   35159: out<=0;
   35160: out<=0;
   35161: out<=1;
   35162: out<=0;
   35163: out<=1;
   35164: out<=0;
   35165: out<=0;
   35166: out<=1;
   35167: out<=1;
   35168: out<=1;
   35169: out<=1;
   35170: out<=0;
   35171: out<=0;
   35172: out<=1;
   35173: out<=0;
   35174: out<=1;
   35175: out<=0;
   35176: out<=0;
   35177: out<=1;
   35178: out<=1;
   35179: out<=0;
   35180: out<=0;
   35181: out<=0;
   35182: out<=0;
   35183: out<=0;
   35184: out<=0;
   35185: out<=1;
   35186: out<=0;
   35187: out<=1;
   35188: out<=1;
   35189: out<=1;
   35190: out<=0;
   35191: out<=0;
   35192: out<=0;
   35193: out<=0;
   35194: out<=0;
   35195: out<=0;
   35196: out<=1;
   35197: out<=0;
   35198: out<=0;
   35199: out<=1;
   35200: out<=0;
   35201: out<=1;
   35202: out<=1;
   35203: out<=0;
   35204: out<=1;
   35205: out<=1;
   35206: out<=1;
   35207: out<=1;
   35208: out<=1;
   35209: out<=1;
   35210: out<=0;
   35211: out<=0;
   35212: out<=0;
   35213: out<=1;
   35214: out<=0;
   35215: out<=1;
   35216: out<=1;
   35217: out<=1;
   35218: out<=1;
   35219: out<=1;
   35220: out<=1;
   35221: out<=0;
   35222: out<=0;
   35223: out<=1;
   35224: out<=1;
   35225: out<=0;
   35226: out<=1;
   35227: out<=0;
   35228: out<=1;
   35229: out<=1;
   35230: out<=0;
   35231: out<=0;
   35232: out<=1;
   35233: out<=1;
   35234: out<=0;
   35235: out<=0;
   35236: out<=1;
   35237: out<=0;
   35238: out<=1;
   35239: out<=0;
   35240: out<=0;
   35241: out<=1;
   35242: out<=1;
   35243: out<=0;
   35244: out<=0;
   35245: out<=0;
   35246: out<=0;
   35247: out<=0;
   35248: out<=0;
   35249: out<=1;
   35250: out<=0;
   35251: out<=1;
   35252: out<=1;
   35253: out<=1;
   35254: out<=0;
   35255: out<=0;
   35256: out<=0;
   35257: out<=0;
   35258: out<=0;
   35259: out<=0;
   35260: out<=1;
   35261: out<=0;
   35262: out<=0;
   35263: out<=1;
   35264: out<=0;
   35265: out<=1;
   35266: out<=1;
   35267: out<=0;
   35268: out<=1;
   35269: out<=1;
   35270: out<=1;
   35271: out<=1;
   35272: out<=1;
   35273: out<=1;
   35274: out<=0;
   35275: out<=0;
   35276: out<=0;
   35277: out<=1;
   35278: out<=0;
   35279: out<=1;
   35280: out<=0;
   35281: out<=0;
   35282: out<=0;
   35283: out<=0;
   35284: out<=0;
   35285: out<=1;
   35286: out<=1;
   35287: out<=0;
   35288: out<=0;
   35289: out<=1;
   35290: out<=0;
   35291: out<=1;
   35292: out<=0;
   35293: out<=0;
   35294: out<=1;
   35295: out<=1;
   35296: out<=0;
   35297: out<=0;
   35298: out<=1;
   35299: out<=1;
   35300: out<=0;
   35301: out<=1;
   35302: out<=0;
   35303: out<=1;
   35304: out<=1;
   35305: out<=0;
   35306: out<=0;
   35307: out<=1;
   35308: out<=1;
   35309: out<=1;
   35310: out<=1;
   35311: out<=1;
   35312: out<=0;
   35313: out<=1;
   35314: out<=0;
   35315: out<=1;
   35316: out<=1;
   35317: out<=1;
   35318: out<=0;
   35319: out<=0;
   35320: out<=0;
   35321: out<=0;
   35322: out<=0;
   35323: out<=0;
   35324: out<=1;
   35325: out<=0;
   35326: out<=0;
   35327: out<=1;
   35328: out<=0;
   35329: out<=1;
   35330: out<=0;
   35331: out<=1;
   35332: out<=1;
   35333: out<=1;
   35334: out<=0;
   35335: out<=0;
   35336: out<=0;
   35337: out<=0;
   35338: out<=0;
   35339: out<=0;
   35340: out<=1;
   35341: out<=0;
   35342: out<=0;
   35343: out<=1;
   35344: out<=0;
   35345: out<=0;
   35346: out<=1;
   35347: out<=1;
   35348: out<=0;
   35349: out<=1;
   35350: out<=0;
   35351: out<=1;
   35352: out<=1;
   35353: out<=0;
   35354: out<=0;
   35355: out<=1;
   35356: out<=1;
   35357: out<=1;
   35358: out<=1;
   35359: out<=1;
   35360: out<=0;
   35361: out<=0;
   35362: out<=0;
   35363: out<=0;
   35364: out<=0;
   35365: out<=1;
   35366: out<=1;
   35367: out<=0;
   35368: out<=0;
   35369: out<=1;
   35370: out<=0;
   35371: out<=1;
   35372: out<=0;
   35373: out<=0;
   35374: out<=1;
   35375: out<=1;
   35376: out<=0;
   35377: out<=1;
   35378: out<=1;
   35379: out<=0;
   35380: out<=1;
   35381: out<=1;
   35382: out<=1;
   35383: out<=1;
   35384: out<=1;
   35385: out<=1;
   35386: out<=0;
   35387: out<=0;
   35388: out<=0;
   35389: out<=1;
   35390: out<=0;
   35391: out<=1;
   35392: out<=0;
   35393: out<=1;
   35394: out<=0;
   35395: out<=1;
   35396: out<=1;
   35397: out<=1;
   35398: out<=0;
   35399: out<=0;
   35400: out<=0;
   35401: out<=0;
   35402: out<=0;
   35403: out<=0;
   35404: out<=1;
   35405: out<=0;
   35406: out<=0;
   35407: out<=1;
   35408: out<=1;
   35409: out<=1;
   35410: out<=0;
   35411: out<=0;
   35412: out<=1;
   35413: out<=0;
   35414: out<=1;
   35415: out<=0;
   35416: out<=0;
   35417: out<=1;
   35418: out<=1;
   35419: out<=0;
   35420: out<=0;
   35421: out<=0;
   35422: out<=0;
   35423: out<=0;
   35424: out<=1;
   35425: out<=1;
   35426: out<=1;
   35427: out<=1;
   35428: out<=1;
   35429: out<=0;
   35430: out<=0;
   35431: out<=1;
   35432: out<=1;
   35433: out<=0;
   35434: out<=1;
   35435: out<=0;
   35436: out<=1;
   35437: out<=1;
   35438: out<=0;
   35439: out<=0;
   35440: out<=0;
   35441: out<=1;
   35442: out<=1;
   35443: out<=0;
   35444: out<=1;
   35445: out<=1;
   35446: out<=1;
   35447: out<=1;
   35448: out<=1;
   35449: out<=1;
   35450: out<=0;
   35451: out<=0;
   35452: out<=0;
   35453: out<=1;
   35454: out<=0;
   35455: out<=1;
   35456: out<=0;
   35457: out<=1;
   35458: out<=0;
   35459: out<=1;
   35460: out<=1;
   35461: out<=1;
   35462: out<=0;
   35463: out<=0;
   35464: out<=0;
   35465: out<=0;
   35466: out<=0;
   35467: out<=0;
   35468: out<=1;
   35469: out<=0;
   35470: out<=0;
   35471: out<=1;
   35472: out<=1;
   35473: out<=1;
   35474: out<=0;
   35475: out<=0;
   35476: out<=1;
   35477: out<=0;
   35478: out<=1;
   35479: out<=0;
   35480: out<=0;
   35481: out<=1;
   35482: out<=1;
   35483: out<=0;
   35484: out<=0;
   35485: out<=0;
   35486: out<=0;
   35487: out<=0;
   35488: out<=0;
   35489: out<=0;
   35490: out<=0;
   35491: out<=0;
   35492: out<=0;
   35493: out<=1;
   35494: out<=1;
   35495: out<=0;
   35496: out<=0;
   35497: out<=1;
   35498: out<=0;
   35499: out<=1;
   35500: out<=0;
   35501: out<=0;
   35502: out<=1;
   35503: out<=1;
   35504: out<=1;
   35505: out<=0;
   35506: out<=0;
   35507: out<=1;
   35508: out<=0;
   35509: out<=0;
   35510: out<=0;
   35511: out<=0;
   35512: out<=0;
   35513: out<=0;
   35514: out<=1;
   35515: out<=1;
   35516: out<=1;
   35517: out<=0;
   35518: out<=1;
   35519: out<=0;
   35520: out<=0;
   35521: out<=1;
   35522: out<=0;
   35523: out<=1;
   35524: out<=1;
   35525: out<=1;
   35526: out<=0;
   35527: out<=0;
   35528: out<=0;
   35529: out<=0;
   35530: out<=0;
   35531: out<=0;
   35532: out<=1;
   35533: out<=0;
   35534: out<=0;
   35535: out<=1;
   35536: out<=0;
   35537: out<=0;
   35538: out<=1;
   35539: out<=1;
   35540: out<=0;
   35541: out<=1;
   35542: out<=0;
   35543: out<=1;
   35544: out<=1;
   35545: out<=0;
   35546: out<=0;
   35547: out<=1;
   35548: out<=1;
   35549: out<=1;
   35550: out<=1;
   35551: out<=1;
   35552: out<=1;
   35553: out<=1;
   35554: out<=1;
   35555: out<=1;
   35556: out<=1;
   35557: out<=0;
   35558: out<=0;
   35559: out<=1;
   35560: out<=1;
   35561: out<=0;
   35562: out<=1;
   35563: out<=0;
   35564: out<=1;
   35565: out<=1;
   35566: out<=0;
   35567: out<=0;
   35568: out<=1;
   35569: out<=0;
   35570: out<=0;
   35571: out<=1;
   35572: out<=0;
   35573: out<=0;
   35574: out<=0;
   35575: out<=0;
   35576: out<=0;
   35577: out<=0;
   35578: out<=1;
   35579: out<=1;
   35580: out<=1;
   35581: out<=0;
   35582: out<=1;
   35583: out<=0;
   35584: out<=1;
   35585: out<=1;
   35586: out<=0;
   35587: out<=0;
   35588: out<=1;
   35589: out<=0;
   35590: out<=1;
   35591: out<=0;
   35592: out<=0;
   35593: out<=1;
   35594: out<=1;
   35595: out<=0;
   35596: out<=0;
   35597: out<=0;
   35598: out<=0;
   35599: out<=0;
   35600: out<=0;
   35601: out<=1;
   35602: out<=0;
   35603: out<=1;
   35604: out<=1;
   35605: out<=1;
   35606: out<=0;
   35607: out<=0;
   35608: out<=0;
   35609: out<=0;
   35610: out<=0;
   35611: out<=0;
   35612: out<=1;
   35613: out<=0;
   35614: out<=0;
   35615: out<=1;
   35616: out<=0;
   35617: out<=1;
   35618: out<=1;
   35619: out<=0;
   35620: out<=1;
   35621: out<=1;
   35622: out<=1;
   35623: out<=1;
   35624: out<=1;
   35625: out<=1;
   35626: out<=0;
   35627: out<=0;
   35628: out<=0;
   35629: out<=1;
   35630: out<=0;
   35631: out<=1;
   35632: out<=1;
   35633: out<=1;
   35634: out<=1;
   35635: out<=1;
   35636: out<=1;
   35637: out<=0;
   35638: out<=0;
   35639: out<=1;
   35640: out<=1;
   35641: out<=0;
   35642: out<=1;
   35643: out<=0;
   35644: out<=1;
   35645: out<=1;
   35646: out<=0;
   35647: out<=0;
   35648: out<=0;
   35649: out<=0;
   35650: out<=1;
   35651: out<=1;
   35652: out<=0;
   35653: out<=1;
   35654: out<=0;
   35655: out<=1;
   35656: out<=1;
   35657: out<=0;
   35658: out<=0;
   35659: out<=1;
   35660: out<=1;
   35661: out<=1;
   35662: out<=1;
   35663: out<=1;
   35664: out<=0;
   35665: out<=1;
   35666: out<=0;
   35667: out<=1;
   35668: out<=1;
   35669: out<=1;
   35670: out<=0;
   35671: out<=0;
   35672: out<=0;
   35673: out<=0;
   35674: out<=0;
   35675: out<=0;
   35676: out<=1;
   35677: out<=0;
   35678: out<=0;
   35679: out<=1;
   35680: out<=0;
   35681: out<=1;
   35682: out<=1;
   35683: out<=0;
   35684: out<=1;
   35685: out<=1;
   35686: out<=1;
   35687: out<=1;
   35688: out<=1;
   35689: out<=1;
   35690: out<=0;
   35691: out<=0;
   35692: out<=0;
   35693: out<=1;
   35694: out<=0;
   35695: out<=1;
   35696: out<=0;
   35697: out<=0;
   35698: out<=0;
   35699: out<=0;
   35700: out<=0;
   35701: out<=1;
   35702: out<=1;
   35703: out<=0;
   35704: out<=0;
   35705: out<=1;
   35706: out<=0;
   35707: out<=1;
   35708: out<=0;
   35709: out<=0;
   35710: out<=1;
   35711: out<=1;
   35712: out<=0;
   35713: out<=0;
   35714: out<=1;
   35715: out<=1;
   35716: out<=0;
   35717: out<=1;
   35718: out<=0;
   35719: out<=1;
   35720: out<=1;
   35721: out<=0;
   35722: out<=0;
   35723: out<=1;
   35724: out<=1;
   35725: out<=1;
   35726: out<=1;
   35727: out<=1;
   35728: out<=0;
   35729: out<=1;
   35730: out<=0;
   35731: out<=1;
   35732: out<=1;
   35733: out<=1;
   35734: out<=0;
   35735: out<=0;
   35736: out<=0;
   35737: out<=0;
   35738: out<=0;
   35739: out<=0;
   35740: out<=1;
   35741: out<=0;
   35742: out<=0;
   35743: out<=1;
   35744: out<=1;
   35745: out<=0;
   35746: out<=0;
   35747: out<=1;
   35748: out<=0;
   35749: out<=0;
   35750: out<=0;
   35751: out<=0;
   35752: out<=0;
   35753: out<=0;
   35754: out<=1;
   35755: out<=1;
   35756: out<=1;
   35757: out<=0;
   35758: out<=1;
   35759: out<=0;
   35760: out<=1;
   35761: out<=1;
   35762: out<=1;
   35763: out<=1;
   35764: out<=1;
   35765: out<=0;
   35766: out<=0;
   35767: out<=1;
   35768: out<=1;
   35769: out<=0;
   35770: out<=1;
   35771: out<=0;
   35772: out<=1;
   35773: out<=1;
   35774: out<=0;
   35775: out<=0;
   35776: out<=1;
   35777: out<=1;
   35778: out<=0;
   35779: out<=0;
   35780: out<=1;
   35781: out<=0;
   35782: out<=1;
   35783: out<=0;
   35784: out<=0;
   35785: out<=1;
   35786: out<=1;
   35787: out<=0;
   35788: out<=0;
   35789: out<=0;
   35790: out<=0;
   35791: out<=0;
   35792: out<=0;
   35793: out<=1;
   35794: out<=0;
   35795: out<=1;
   35796: out<=1;
   35797: out<=1;
   35798: out<=0;
   35799: out<=0;
   35800: out<=0;
   35801: out<=0;
   35802: out<=0;
   35803: out<=0;
   35804: out<=1;
   35805: out<=0;
   35806: out<=0;
   35807: out<=1;
   35808: out<=1;
   35809: out<=0;
   35810: out<=0;
   35811: out<=1;
   35812: out<=0;
   35813: out<=0;
   35814: out<=0;
   35815: out<=0;
   35816: out<=0;
   35817: out<=0;
   35818: out<=1;
   35819: out<=1;
   35820: out<=1;
   35821: out<=0;
   35822: out<=1;
   35823: out<=0;
   35824: out<=0;
   35825: out<=0;
   35826: out<=0;
   35827: out<=0;
   35828: out<=0;
   35829: out<=1;
   35830: out<=1;
   35831: out<=0;
   35832: out<=0;
   35833: out<=1;
   35834: out<=0;
   35835: out<=1;
   35836: out<=0;
   35837: out<=0;
   35838: out<=1;
   35839: out<=1;
   35840: out<=0;
   35841: out<=1;
   35842: out<=1;
   35843: out<=0;
   35844: out<=0;
   35845: out<=0;
   35846: out<=0;
   35847: out<=0;
   35848: out<=0;
   35849: out<=0;
   35850: out<=1;
   35851: out<=1;
   35852: out<=0;
   35853: out<=1;
   35854: out<=0;
   35855: out<=1;
   35856: out<=1;
   35857: out<=1;
   35858: out<=1;
   35859: out<=1;
   35860: out<=0;
   35861: out<=1;
   35862: out<=1;
   35863: out<=0;
   35864: out<=0;
   35865: out<=1;
   35866: out<=0;
   35867: out<=1;
   35868: out<=1;
   35869: out<=1;
   35870: out<=0;
   35871: out<=0;
   35872: out<=0;
   35873: out<=0;
   35874: out<=1;
   35875: out<=1;
   35876: out<=1;
   35877: out<=0;
   35878: out<=1;
   35879: out<=0;
   35880: out<=0;
   35881: out<=1;
   35882: out<=1;
   35883: out<=0;
   35884: out<=1;
   35885: out<=1;
   35886: out<=1;
   35887: out<=1;
   35888: out<=1;
   35889: out<=0;
   35890: out<=1;
   35891: out<=0;
   35892: out<=1;
   35893: out<=1;
   35894: out<=0;
   35895: out<=0;
   35896: out<=0;
   35897: out<=0;
   35898: out<=0;
   35899: out<=0;
   35900: out<=0;
   35901: out<=1;
   35902: out<=1;
   35903: out<=0;
   35904: out<=0;
   35905: out<=1;
   35906: out<=1;
   35907: out<=0;
   35908: out<=0;
   35909: out<=0;
   35910: out<=0;
   35911: out<=0;
   35912: out<=0;
   35913: out<=0;
   35914: out<=1;
   35915: out<=1;
   35916: out<=0;
   35917: out<=1;
   35918: out<=0;
   35919: out<=1;
   35920: out<=0;
   35921: out<=0;
   35922: out<=0;
   35923: out<=0;
   35924: out<=1;
   35925: out<=0;
   35926: out<=0;
   35927: out<=1;
   35928: out<=1;
   35929: out<=0;
   35930: out<=1;
   35931: out<=0;
   35932: out<=0;
   35933: out<=0;
   35934: out<=1;
   35935: out<=1;
   35936: out<=1;
   35937: out<=1;
   35938: out<=0;
   35939: out<=0;
   35940: out<=0;
   35941: out<=1;
   35942: out<=0;
   35943: out<=1;
   35944: out<=1;
   35945: out<=0;
   35946: out<=0;
   35947: out<=1;
   35948: out<=0;
   35949: out<=0;
   35950: out<=0;
   35951: out<=0;
   35952: out<=1;
   35953: out<=0;
   35954: out<=1;
   35955: out<=0;
   35956: out<=1;
   35957: out<=1;
   35958: out<=0;
   35959: out<=0;
   35960: out<=0;
   35961: out<=0;
   35962: out<=0;
   35963: out<=0;
   35964: out<=0;
   35965: out<=1;
   35966: out<=1;
   35967: out<=0;
   35968: out<=1;
   35969: out<=0;
   35970: out<=0;
   35971: out<=1;
   35972: out<=1;
   35973: out<=1;
   35974: out<=1;
   35975: out<=1;
   35976: out<=1;
   35977: out<=1;
   35978: out<=0;
   35979: out<=0;
   35980: out<=1;
   35981: out<=0;
   35982: out<=1;
   35983: out<=0;
   35984: out<=1;
   35985: out<=1;
   35986: out<=1;
   35987: out<=1;
   35988: out<=0;
   35989: out<=1;
   35990: out<=1;
   35991: out<=0;
   35992: out<=0;
   35993: out<=1;
   35994: out<=0;
   35995: out<=1;
   35996: out<=1;
   35997: out<=1;
   35998: out<=0;
   35999: out<=0;
   36000: out<=1;
   36001: out<=1;
   36002: out<=0;
   36003: out<=0;
   36004: out<=0;
   36005: out<=1;
   36006: out<=0;
   36007: out<=1;
   36008: out<=1;
   36009: out<=0;
   36010: out<=0;
   36011: out<=1;
   36012: out<=0;
   36013: out<=0;
   36014: out<=0;
   36015: out<=0;
   36016: out<=1;
   36017: out<=0;
   36018: out<=1;
   36019: out<=0;
   36020: out<=1;
   36021: out<=1;
   36022: out<=0;
   36023: out<=0;
   36024: out<=0;
   36025: out<=0;
   36026: out<=0;
   36027: out<=0;
   36028: out<=0;
   36029: out<=1;
   36030: out<=1;
   36031: out<=0;
   36032: out<=1;
   36033: out<=0;
   36034: out<=0;
   36035: out<=1;
   36036: out<=1;
   36037: out<=1;
   36038: out<=1;
   36039: out<=1;
   36040: out<=1;
   36041: out<=1;
   36042: out<=0;
   36043: out<=0;
   36044: out<=1;
   36045: out<=0;
   36046: out<=1;
   36047: out<=0;
   36048: out<=0;
   36049: out<=0;
   36050: out<=0;
   36051: out<=0;
   36052: out<=1;
   36053: out<=0;
   36054: out<=0;
   36055: out<=1;
   36056: out<=1;
   36057: out<=0;
   36058: out<=1;
   36059: out<=0;
   36060: out<=0;
   36061: out<=0;
   36062: out<=1;
   36063: out<=1;
   36064: out<=0;
   36065: out<=0;
   36066: out<=1;
   36067: out<=1;
   36068: out<=1;
   36069: out<=0;
   36070: out<=1;
   36071: out<=0;
   36072: out<=0;
   36073: out<=1;
   36074: out<=1;
   36075: out<=0;
   36076: out<=1;
   36077: out<=1;
   36078: out<=1;
   36079: out<=1;
   36080: out<=1;
   36081: out<=0;
   36082: out<=1;
   36083: out<=0;
   36084: out<=1;
   36085: out<=1;
   36086: out<=0;
   36087: out<=0;
   36088: out<=0;
   36089: out<=0;
   36090: out<=0;
   36091: out<=0;
   36092: out<=0;
   36093: out<=1;
   36094: out<=1;
   36095: out<=0;
   36096: out<=0;
   36097: out<=0;
   36098: out<=0;
   36099: out<=0;
   36100: out<=1;
   36101: out<=0;
   36102: out<=0;
   36103: out<=1;
   36104: out<=1;
   36105: out<=0;
   36106: out<=1;
   36107: out<=0;
   36108: out<=0;
   36109: out<=0;
   36110: out<=1;
   36111: out<=1;
   36112: out<=0;
   36113: out<=1;
   36114: out<=1;
   36115: out<=0;
   36116: out<=0;
   36117: out<=0;
   36118: out<=0;
   36119: out<=0;
   36120: out<=0;
   36121: out<=0;
   36122: out<=1;
   36123: out<=1;
   36124: out<=0;
   36125: out<=1;
   36126: out<=0;
   36127: out<=1;
   36128: out<=1;
   36129: out<=0;
   36130: out<=1;
   36131: out<=0;
   36132: out<=1;
   36133: out<=1;
   36134: out<=0;
   36135: out<=0;
   36136: out<=0;
   36137: out<=0;
   36138: out<=0;
   36139: out<=0;
   36140: out<=0;
   36141: out<=1;
   36142: out<=1;
   36143: out<=0;
   36144: out<=1;
   36145: out<=1;
   36146: out<=0;
   36147: out<=0;
   36148: out<=0;
   36149: out<=1;
   36150: out<=0;
   36151: out<=1;
   36152: out<=1;
   36153: out<=0;
   36154: out<=0;
   36155: out<=1;
   36156: out<=0;
   36157: out<=0;
   36158: out<=0;
   36159: out<=0;
   36160: out<=1;
   36161: out<=1;
   36162: out<=1;
   36163: out<=1;
   36164: out<=0;
   36165: out<=1;
   36166: out<=1;
   36167: out<=0;
   36168: out<=0;
   36169: out<=1;
   36170: out<=0;
   36171: out<=1;
   36172: out<=1;
   36173: out<=1;
   36174: out<=0;
   36175: out<=0;
   36176: out<=0;
   36177: out<=1;
   36178: out<=1;
   36179: out<=0;
   36180: out<=0;
   36181: out<=0;
   36182: out<=0;
   36183: out<=0;
   36184: out<=0;
   36185: out<=0;
   36186: out<=1;
   36187: out<=1;
   36188: out<=0;
   36189: out<=1;
   36190: out<=0;
   36191: out<=1;
   36192: out<=1;
   36193: out<=0;
   36194: out<=1;
   36195: out<=0;
   36196: out<=1;
   36197: out<=1;
   36198: out<=0;
   36199: out<=0;
   36200: out<=0;
   36201: out<=0;
   36202: out<=0;
   36203: out<=0;
   36204: out<=0;
   36205: out<=1;
   36206: out<=1;
   36207: out<=0;
   36208: out<=0;
   36209: out<=0;
   36210: out<=1;
   36211: out<=1;
   36212: out<=1;
   36213: out<=0;
   36214: out<=1;
   36215: out<=0;
   36216: out<=0;
   36217: out<=1;
   36218: out<=1;
   36219: out<=0;
   36220: out<=1;
   36221: out<=1;
   36222: out<=1;
   36223: out<=1;
   36224: out<=0;
   36225: out<=0;
   36226: out<=0;
   36227: out<=0;
   36228: out<=1;
   36229: out<=0;
   36230: out<=0;
   36231: out<=1;
   36232: out<=1;
   36233: out<=0;
   36234: out<=1;
   36235: out<=0;
   36236: out<=0;
   36237: out<=0;
   36238: out<=1;
   36239: out<=1;
   36240: out<=1;
   36241: out<=0;
   36242: out<=0;
   36243: out<=1;
   36244: out<=1;
   36245: out<=1;
   36246: out<=1;
   36247: out<=1;
   36248: out<=1;
   36249: out<=1;
   36250: out<=0;
   36251: out<=0;
   36252: out<=1;
   36253: out<=0;
   36254: out<=1;
   36255: out<=0;
   36256: out<=1;
   36257: out<=0;
   36258: out<=1;
   36259: out<=0;
   36260: out<=1;
   36261: out<=1;
   36262: out<=0;
   36263: out<=0;
   36264: out<=0;
   36265: out<=0;
   36266: out<=0;
   36267: out<=0;
   36268: out<=0;
   36269: out<=1;
   36270: out<=1;
   36271: out<=0;
   36272: out<=0;
   36273: out<=0;
   36274: out<=1;
   36275: out<=1;
   36276: out<=1;
   36277: out<=0;
   36278: out<=1;
   36279: out<=0;
   36280: out<=0;
   36281: out<=1;
   36282: out<=1;
   36283: out<=0;
   36284: out<=1;
   36285: out<=1;
   36286: out<=1;
   36287: out<=1;
   36288: out<=1;
   36289: out<=1;
   36290: out<=1;
   36291: out<=1;
   36292: out<=0;
   36293: out<=1;
   36294: out<=1;
   36295: out<=0;
   36296: out<=0;
   36297: out<=1;
   36298: out<=0;
   36299: out<=1;
   36300: out<=1;
   36301: out<=1;
   36302: out<=0;
   36303: out<=0;
   36304: out<=1;
   36305: out<=0;
   36306: out<=0;
   36307: out<=1;
   36308: out<=1;
   36309: out<=1;
   36310: out<=1;
   36311: out<=1;
   36312: out<=1;
   36313: out<=1;
   36314: out<=0;
   36315: out<=0;
   36316: out<=1;
   36317: out<=0;
   36318: out<=1;
   36319: out<=0;
   36320: out<=1;
   36321: out<=0;
   36322: out<=1;
   36323: out<=0;
   36324: out<=1;
   36325: out<=1;
   36326: out<=0;
   36327: out<=0;
   36328: out<=0;
   36329: out<=0;
   36330: out<=0;
   36331: out<=0;
   36332: out<=0;
   36333: out<=1;
   36334: out<=1;
   36335: out<=0;
   36336: out<=1;
   36337: out<=1;
   36338: out<=0;
   36339: out<=0;
   36340: out<=0;
   36341: out<=1;
   36342: out<=0;
   36343: out<=1;
   36344: out<=1;
   36345: out<=0;
   36346: out<=0;
   36347: out<=1;
   36348: out<=0;
   36349: out<=0;
   36350: out<=0;
   36351: out<=0;
   36352: out<=1;
   36353: out<=1;
   36354: out<=0;
   36355: out<=0;
   36356: out<=0;
   36357: out<=1;
   36358: out<=0;
   36359: out<=1;
   36360: out<=1;
   36361: out<=0;
   36362: out<=0;
   36363: out<=1;
   36364: out<=0;
   36365: out<=0;
   36366: out<=0;
   36367: out<=0;
   36368: out<=1;
   36369: out<=0;
   36370: out<=1;
   36371: out<=0;
   36372: out<=1;
   36373: out<=1;
   36374: out<=0;
   36375: out<=0;
   36376: out<=0;
   36377: out<=0;
   36378: out<=0;
   36379: out<=0;
   36380: out<=0;
   36381: out<=1;
   36382: out<=1;
   36383: out<=0;
   36384: out<=1;
   36385: out<=0;
   36386: out<=0;
   36387: out<=1;
   36388: out<=1;
   36389: out<=1;
   36390: out<=1;
   36391: out<=1;
   36392: out<=1;
   36393: out<=1;
   36394: out<=0;
   36395: out<=0;
   36396: out<=1;
   36397: out<=0;
   36398: out<=1;
   36399: out<=0;
   36400: out<=1;
   36401: out<=1;
   36402: out<=1;
   36403: out<=1;
   36404: out<=0;
   36405: out<=1;
   36406: out<=1;
   36407: out<=0;
   36408: out<=0;
   36409: out<=1;
   36410: out<=0;
   36411: out<=1;
   36412: out<=1;
   36413: out<=1;
   36414: out<=0;
   36415: out<=0;
   36416: out<=0;
   36417: out<=0;
   36418: out<=1;
   36419: out<=1;
   36420: out<=1;
   36421: out<=0;
   36422: out<=1;
   36423: out<=0;
   36424: out<=0;
   36425: out<=1;
   36426: out<=1;
   36427: out<=0;
   36428: out<=1;
   36429: out<=1;
   36430: out<=1;
   36431: out<=1;
   36432: out<=1;
   36433: out<=0;
   36434: out<=1;
   36435: out<=0;
   36436: out<=1;
   36437: out<=1;
   36438: out<=0;
   36439: out<=0;
   36440: out<=0;
   36441: out<=0;
   36442: out<=0;
   36443: out<=0;
   36444: out<=0;
   36445: out<=1;
   36446: out<=1;
   36447: out<=0;
   36448: out<=1;
   36449: out<=0;
   36450: out<=0;
   36451: out<=1;
   36452: out<=1;
   36453: out<=1;
   36454: out<=1;
   36455: out<=1;
   36456: out<=1;
   36457: out<=1;
   36458: out<=0;
   36459: out<=0;
   36460: out<=1;
   36461: out<=0;
   36462: out<=1;
   36463: out<=0;
   36464: out<=0;
   36465: out<=0;
   36466: out<=0;
   36467: out<=0;
   36468: out<=1;
   36469: out<=0;
   36470: out<=0;
   36471: out<=1;
   36472: out<=1;
   36473: out<=0;
   36474: out<=1;
   36475: out<=0;
   36476: out<=0;
   36477: out<=0;
   36478: out<=1;
   36479: out<=1;
   36480: out<=0;
   36481: out<=0;
   36482: out<=1;
   36483: out<=1;
   36484: out<=1;
   36485: out<=0;
   36486: out<=1;
   36487: out<=0;
   36488: out<=0;
   36489: out<=1;
   36490: out<=1;
   36491: out<=0;
   36492: out<=1;
   36493: out<=1;
   36494: out<=1;
   36495: out<=1;
   36496: out<=1;
   36497: out<=0;
   36498: out<=1;
   36499: out<=0;
   36500: out<=1;
   36501: out<=1;
   36502: out<=0;
   36503: out<=0;
   36504: out<=0;
   36505: out<=0;
   36506: out<=0;
   36507: out<=0;
   36508: out<=0;
   36509: out<=1;
   36510: out<=1;
   36511: out<=0;
   36512: out<=0;
   36513: out<=1;
   36514: out<=1;
   36515: out<=0;
   36516: out<=0;
   36517: out<=0;
   36518: out<=0;
   36519: out<=0;
   36520: out<=0;
   36521: out<=0;
   36522: out<=1;
   36523: out<=1;
   36524: out<=0;
   36525: out<=1;
   36526: out<=0;
   36527: out<=1;
   36528: out<=1;
   36529: out<=1;
   36530: out<=1;
   36531: out<=1;
   36532: out<=0;
   36533: out<=1;
   36534: out<=1;
   36535: out<=0;
   36536: out<=0;
   36537: out<=1;
   36538: out<=0;
   36539: out<=1;
   36540: out<=1;
   36541: out<=1;
   36542: out<=0;
   36543: out<=0;
   36544: out<=1;
   36545: out<=1;
   36546: out<=0;
   36547: out<=0;
   36548: out<=0;
   36549: out<=1;
   36550: out<=0;
   36551: out<=1;
   36552: out<=1;
   36553: out<=0;
   36554: out<=0;
   36555: out<=1;
   36556: out<=0;
   36557: out<=0;
   36558: out<=0;
   36559: out<=0;
   36560: out<=1;
   36561: out<=0;
   36562: out<=1;
   36563: out<=0;
   36564: out<=1;
   36565: out<=1;
   36566: out<=0;
   36567: out<=0;
   36568: out<=0;
   36569: out<=0;
   36570: out<=0;
   36571: out<=0;
   36572: out<=0;
   36573: out<=1;
   36574: out<=1;
   36575: out<=0;
   36576: out<=0;
   36577: out<=1;
   36578: out<=1;
   36579: out<=0;
   36580: out<=0;
   36581: out<=0;
   36582: out<=0;
   36583: out<=0;
   36584: out<=0;
   36585: out<=0;
   36586: out<=1;
   36587: out<=1;
   36588: out<=0;
   36589: out<=1;
   36590: out<=0;
   36591: out<=1;
   36592: out<=0;
   36593: out<=0;
   36594: out<=0;
   36595: out<=0;
   36596: out<=1;
   36597: out<=0;
   36598: out<=0;
   36599: out<=1;
   36600: out<=1;
   36601: out<=0;
   36602: out<=1;
   36603: out<=0;
   36604: out<=0;
   36605: out<=0;
   36606: out<=1;
   36607: out<=1;
   36608: out<=1;
   36609: out<=0;
   36610: out<=1;
   36611: out<=0;
   36612: out<=1;
   36613: out<=1;
   36614: out<=0;
   36615: out<=0;
   36616: out<=0;
   36617: out<=0;
   36618: out<=0;
   36619: out<=0;
   36620: out<=0;
   36621: out<=1;
   36622: out<=1;
   36623: out<=0;
   36624: out<=0;
   36625: out<=0;
   36626: out<=1;
   36627: out<=1;
   36628: out<=1;
   36629: out<=0;
   36630: out<=1;
   36631: out<=0;
   36632: out<=0;
   36633: out<=1;
   36634: out<=1;
   36635: out<=0;
   36636: out<=1;
   36637: out<=1;
   36638: out<=1;
   36639: out<=1;
   36640: out<=0;
   36641: out<=0;
   36642: out<=0;
   36643: out<=0;
   36644: out<=1;
   36645: out<=0;
   36646: out<=0;
   36647: out<=1;
   36648: out<=1;
   36649: out<=0;
   36650: out<=1;
   36651: out<=0;
   36652: out<=0;
   36653: out<=0;
   36654: out<=1;
   36655: out<=1;
   36656: out<=1;
   36657: out<=0;
   36658: out<=0;
   36659: out<=1;
   36660: out<=1;
   36661: out<=1;
   36662: out<=1;
   36663: out<=1;
   36664: out<=1;
   36665: out<=1;
   36666: out<=0;
   36667: out<=0;
   36668: out<=1;
   36669: out<=0;
   36670: out<=1;
   36671: out<=0;
   36672: out<=1;
   36673: out<=0;
   36674: out<=1;
   36675: out<=0;
   36676: out<=1;
   36677: out<=1;
   36678: out<=0;
   36679: out<=0;
   36680: out<=0;
   36681: out<=0;
   36682: out<=0;
   36683: out<=0;
   36684: out<=0;
   36685: out<=1;
   36686: out<=1;
   36687: out<=0;
   36688: out<=1;
   36689: out<=1;
   36690: out<=0;
   36691: out<=0;
   36692: out<=0;
   36693: out<=1;
   36694: out<=0;
   36695: out<=1;
   36696: out<=1;
   36697: out<=0;
   36698: out<=0;
   36699: out<=1;
   36700: out<=0;
   36701: out<=0;
   36702: out<=0;
   36703: out<=0;
   36704: out<=1;
   36705: out<=1;
   36706: out<=1;
   36707: out<=1;
   36708: out<=0;
   36709: out<=1;
   36710: out<=1;
   36711: out<=0;
   36712: out<=0;
   36713: out<=1;
   36714: out<=0;
   36715: out<=1;
   36716: out<=1;
   36717: out<=1;
   36718: out<=0;
   36719: out<=0;
   36720: out<=1;
   36721: out<=0;
   36722: out<=0;
   36723: out<=1;
   36724: out<=1;
   36725: out<=1;
   36726: out<=1;
   36727: out<=1;
   36728: out<=1;
   36729: out<=1;
   36730: out<=0;
   36731: out<=0;
   36732: out<=1;
   36733: out<=0;
   36734: out<=1;
   36735: out<=0;
   36736: out<=1;
   36737: out<=0;
   36738: out<=1;
   36739: out<=0;
   36740: out<=1;
   36741: out<=1;
   36742: out<=0;
   36743: out<=0;
   36744: out<=0;
   36745: out<=0;
   36746: out<=0;
   36747: out<=0;
   36748: out<=0;
   36749: out<=1;
   36750: out<=1;
   36751: out<=0;
   36752: out<=1;
   36753: out<=1;
   36754: out<=0;
   36755: out<=0;
   36756: out<=0;
   36757: out<=1;
   36758: out<=0;
   36759: out<=1;
   36760: out<=1;
   36761: out<=0;
   36762: out<=0;
   36763: out<=1;
   36764: out<=0;
   36765: out<=0;
   36766: out<=0;
   36767: out<=0;
   36768: out<=0;
   36769: out<=0;
   36770: out<=0;
   36771: out<=0;
   36772: out<=1;
   36773: out<=0;
   36774: out<=0;
   36775: out<=1;
   36776: out<=1;
   36777: out<=0;
   36778: out<=1;
   36779: out<=0;
   36780: out<=0;
   36781: out<=0;
   36782: out<=1;
   36783: out<=1;
   36784: out<=0;
   36785: out<=1;
   36786: out<=1;
   36787: out<=0;
   36788: out<=0;
   36789: out<=0;
   36790: out<=0;
   36791: out<=0;
   36792: out<=0;
   36793: out<=0;
   36794: out<=1;
   36795: out<=1;
   36796: out<=0;
   36797: out<=1;
   36798: out<=0;
   36799: out<=1;
   36800: out<=1;
   36801: out<=0;
   36802: out<=1;
   36803: out<=0;
   36804: out<=1;
   36805: out<=1;
   36806: out<=0;
   36807: out<=0;
   36808: out<=0;
   36809: out<=0;
   36810: out<=0;
   36811: out<=0;
   36812: out<=0;
   36813: out<=1;
   36814: out<=1;
   36815: out<=0;
   36816: out<=0;
   36817: out<=0;
   36818: out<=1;
   36819: out<=1;
   36820: out<=1;
   36821: out<=0;
   36822: out<=1;
   36823: out<=0;
   36824: out<=0;
   36825: out<=1;
   36826: out<=1;
   36827: out<=0;
   36828: out<=1;
   36829: out<=1;
   36830: out<=1;
   36831: out<=1;
   36832: out<=1;
   36833: out<=1;
   36834: out<=1;
   36835: out<=1;
   36836: out<=0;
   36837: out<=1;
   36838: out<=1;
   36839: out<=0;
   36840: out<=0;
   36841: out<=1;
   36842: out<=0;
   36843: out<=1;
   36844: out<=1;
   36845: out<=1;
   36846: out<=0;
   36847: out<=0;
   36848: out<=0;
   36849: out<=1;
   36850: out<=1;
   36851: out<=0;
   36852: out<=0;
   36853: out<=0;
   36854: out<=0;
   36855: out<=0;
   36856: out<=0;
   36857: out<=0;
   36858: out<=1;
   36859: out<=1;
   36860: out<=0;
   36861: out<=1;
   36862: out<=0;
   36863: out<=1;
   36864: out<=0;
   36865: out<=1;
   36866: out<=0;
   36867: out<=1;
   36868: out<=1;
   36869: out<=1;
   36870: out<=0;
   36871: out<=0;
   36872: out<=1;
   36873: out<=1;
   36874: out<=1;
   36875: out<=1;
   36876: out<=0;
   36877: out<=1;
   36878: out<=1;
   36879: out<=0;
   36880: out<=1;
   36881: out<=1;
   36882: out<=0;
   36883: out<=0;
   36884: out<=1;
   36885: out<=0;
   36886: out<=1;
   36887: out<=0;
   36888: out<=1;
   36889: out<=0;
   36890: out<=0;
   36891: out<=1;
   36892: out<=1;
   36893: out<=1;
   36894: out<=1;
   36895: out<=1;
   36896: out<=0;
   36897: out<=0;
   36898: out<=0;
   36899: out<=0;
   36900: out<=0;
   36901: out<=1;
   36902: out<=1;
   36903: out<=0;
   36904: out<=1;
   36905: out<=0;
   36906: out<=1;
   36907: out<=0;
   36908: out<=1;
   36909: out<=1;
   36910: out<=0;
   36911: out<=0;
   36912: out<=1;
   36913: out<=0;
   36914: out<=0;
   36915: out<=1;
   36916: out<=0;
   36917: out<=0;
   36918: out<=0;
   36919: out<=0;
   36920: out<=1;
   36921: out<=1;
   36922: out<=0;
   36923: out<=0;
   36924: out<=0;
   36925: out<=1;
   36926: out<=0;
   36927: out<=1;
   36928: out<=0;
   36929: out<=1;
   36930: out<=0;
   36931: out<=1;
   36932: out<=1;
   36933: out<=1;
   36934: out<=0;
   36935: out<=0;
   36936: out<=1;
   36937: out<=1;
   36938: out<=1;
   36939: out<=1;
   36940: out<=0;
   36941: out<=1;
   36942: out<=1;
   36943: out<=0;
   36944: out<=0;
   36945: out<=0;
   36946: out<=1;
   36947: out<=1;
   36948: out<=0;
   36949: out<=1;
   36950: out<=0;
   36951: out<=1;
   36952: out<=0;
   36953: out<=1;
   36954: out<=1;
   36955: out<=0;
   36956: out<=0;
   36957: out<=0;
   36958: out<=0;
   36959: out<=0;
   36960: out<=1;
   36961: out<=1;
   36962: out<=1;
   36963: out<=1;
   36964: out<=1;
   36965: out<=0;
   36966: out<=0;
   36967: out<=1;
   36968: out<=0;
   36969: out<=1;
   36970: out<=0;
   36971: out<=1;
   36972: out<=0;
   36973: out<=0;
   36974: out<=1;
   36975: out<=1;
   36976: out<=1;
   36977: out<=0;
   36978: out<=0;
   36979: out<=1;
   36980: out<=0;
   36981: out<=0;
   36982: out<=0;
   36983: out<=0;
   36984: out<=1;
   36985: out<=1;
   36986: out<=0;
   36987: out<=0;
   36988: out<=0;
   36989: out<=1;
   36990: out<=0;
   36991: out<=1;
   36992: out<=0;
   36993: out<=1;
   36994: out<=0;
   36995: out<=1;
   36996: out<=1;
   36997: out<=1;
   36998: out<=0;
   36999: out<=0;
   37000: out<=1;
   37001: out<=1;
   37002: out<=1;
   37003: out<=1;
   37004: out<=0;
   37005: out<=1;
   37006: out<=1;
   37007: out<=0;
   37008: out<=0;
   37009: out<=0;
   37010: out<=1;
   37011: out<=1;
   37012: out<=0;
   37013: out<=1;
   37014: out<=0;
   37015: out<=1;
   37016: out<=0;
   37017: out<=1;
   37018: out<=1;
   37019: out<=0;
   37020: out<=0;
   37021: out<=0;
   37022: out<=0;
   37023: out<=0;
   37024: out<=0;
   37025: out<=0;
   37026: out<=0;
   37027: out<=0;
   37028: out<=0;
   37029: out<=1;
   37030: out<=1;
   37031: out<=0;
   37032: out<=1;
   37033: out<=0;
   37034: out<=1;
   37035: out<=0;
   37036: out<=1;
   37037: out<=1;
   37038: out<=0;
   37039: out<=0;
   37040: out<=0;
   37041: out<=1;
   37042: out<=1;
   37043: out<=0;
   37044: out<=1;
   37045: out<=1;
   37046: out<=1;
   37047: out<=1;
   37048: out<=0;
   37049: out<=0;
   37050: out<=1;
   37051: out<=1;
   37052: out<=1;
   37053: out<=0;
   37054: out<=1;
   37055: out<=0;
   37056: out<=0;
   37057: out<=1;
   37058: out<=0;
   37059: out<=1;
   37060: out<=1;
   37061: out<=1;
   37062: out<=0;
   37063: out<=0;
   37064: out<=1;
   37065: out<=1;
   37066: out<=1;
   37067: out<=1;
   37068: out<=0;
   37069: out<=1;
   37070: out<=1;
   37071: out<=0;
   37072: out<=1;
   37073: out<=1;
   37074: out<=0;
   37075: out<=0;
   37076: out<=1;
   37077: out<=0;
   37078: out<=1;
   37079: out<=0;
   37080: out<=1;
   37081: out<=0;
   37082: out<=0;
   37083: out<=1;
   37084: out<=1;
   37085: out<=1;
   37086: out<=1;
   37087: out<=1;
   37088: out<=1;
   37089: out<=1;
   37090: out<=1;
   37091: out<=1;
   37092: out<=1;
   37093: out<=0;
   37094: out<=0;
   37095: out<=1;
   37096: out<=0;
   37097: out<=1;
   37098: out<=0;
   37099: out<=1;
   37100: out<=0;
   37101: out<=0;
   37102: out<=1;
   37103: out<=1;
   37104: out<=0;
   37105: out<=1;
   37106: out<=1;
   37107: out<=0;
   37108: out<=1;
   37109: out<=1;
   37110: out<=1;
   37111: out<=1;
   37112: out<=0;
   37113: out<=0;
   37114: out<=1;
   37115: out<=1;
   37116: out<=1;
   37117: out<=0;
   37118: out<=1;
   37119: out<=0;
   37120: out<=0;
   37121: out<=0;
   37122: out<=1;
   37123: out<=1;
   37124: out<=0;
   37125: out<=1;
   37126: out<=0;
   37127: out<=1;
   37128: out<=0;
   37129: out<=1;
   37130: out<=1;
   37131: out<=0;
   37132: out<=0;
   37133: out<=0;
   37134: out<=0;
   37135: out<=0;
   37136: out<=0;
   37137: out<=1;
   37138: out<=0;
   37139: out<=1;
   37140: out<=1;
   37141: out<=1;
   37142: out<=0;
   37143: out<=0;
   37144: out<=1;
   37145: out<=1;
   37146: out<=1;
   37147: out<=1;
   37148: out<=0;
   37149: out<=1;
   37150: out<=1;
   37151: out<=0;
   37152: out<=1;
   37153: out<=0;
   37154: out<=0;
   37155: out<=1;
   37156: out<=0;
   37157: out<=0;
   37158: out<=0;
   37159: out<=0;
   37160: out<=1;
   37161: out<=1;
   37162: out<=0;
   37163: out<=0;
   37164: out<=0;
   37165: out<=1;
   37166: out<=0;
   37167: out<=1;
   37168: out<=1;
   37169: out<=1;
   37170: out<=1;
   37171: out<=1;
   37172: out<=1;
   37173: out<=0;
   37174: out<=0;
   37175: out<=1;
   37176: out<=0;
   37177: out<=1;
   37178: out<=0;
   37179: out<=1;
   37180: out<=0;
   37181: out<=0;
   37182: out<=1;
   37183: out<=1;
   37184: out<=1;
   37185: out<=1;
   37186: out<=0;
   37187: out<=0;
   37188: out<=1;
   37189: out<=0;
   37190: out<=1;
   37191: out<=0;
   37192: out<=1;
   37193: out<=0;
   37194: out<=0;
   37195: out<=1;
   37196: out<=1;
   37197: out<=1;
   37198: out<=1;
   37199: out<=1;
   37200: out<=0;
   37201: out<=1;
   37202: out<=0;
   37203: out<=1;
   37204: out<=1;
   37205: out<=1;
   37206: out<=0;
   37207: out<=0;
   37208: out<=1;
   37209: out<=1;
   37210: out<=1;
   37211: out<=1;
   37212: out<=0;
   37213: out<=1;
   37214: out<=1;
   37215: out<=0;
   37216: out<=1;
   37217: out<=0;
   37218: out<=0;
   37219: out<=1;
   37220: out<=0;
   37221: out<=0;
   37222: out<=0;
   37223: out<=0;
   37224: out<=1;
   37225: out<=1;
   37226: out<=0;
   37227: out<=0;
   37228: out<=0;
   37229: out<=1;
   37230: out<=0;
   37231: out<=1;
   37232: out<=0;
   37233: out<=0;
   37234: out<=0;
   37235: out<=0;
   37236: out<=0;
   37237: out<=1;
   37238: out<=1;
   37239: out<=0;
   37240: out<=1;
   37241: out<=0;
   37242: out<=1;
   37243: out<=0;
   37244: out<=1;
   37245: out<=1;
   37246: out<=0;
   37247: out<=0;
   37248: out<=1;
   37249: out<=1;
   37250: out<=0;
   37251: out<=0;
   37252: out<=1;
   37253: out<=0;
   37254: out<=1;
   37255: out<=0;
   37256: out<=1;
   37257: out<=0;
   37258: out<=0;
   37259: out<=1;
   37260: out<=1;
   37261: out<=1;
   37262: out<=1;
   37263: out<=1;
   37264: out<=0;
   37265: out<=1;
   37266: out<=0;
   37267: out<=1;
   37268: out<=1;
   37269: out<=1;
   37270: out<=0;
   37271: out<=0;
   37272: out<=1;
   37273: out<=1;
   37274: out<=1;
   37275: out<=1;
   37276: out<=0;
   37277: out<=1;
   37278: out<=1;
   37279: out<=0;
   37280: out<=0;
   37281: out<=1;
   37282: out<=1;
   37283: out<=0;
   37284: out<=1;
   37285: out<=1;
   37286: out<=1;
   37287: out<=1;
   37288: out<=0;
   37289: out<=0;
   37290: out<=1;
   37291: out<=1;
   37292: out<=1;
   37293: out<=0;
   37294: out<=1;
   37295: out<=0;
   37296: out<=1;
   37297: out<=1;
   37298: out<=1;
   37299: out<=1;
   37300: out<=1;
   37301: out<=0;
   37302: out<=0;
   37303: out<=1;
   37304: out<=0;
   37305: out<=1;
   37306: out<=0;
   37307: out<=1;
   37308: out<=0;
   37309: out<=0;
   37310: out<=1;
   37311: out<=1;
   37312: out<=0;
   37313: out<=0;
   37314: out<=1;
   37315: out<=1;
   37316: out<=0;
   37317: out<=1;
   37318: out<=0;
   37319: out<=1;
   37320: out<=0;
   37321: out<=1;
   37322: out<=1;
   37323: out<=0;
   37324: out<=0;
   37325: out<=0;
   37326: out<=0;
   37327: out<=0;
   37328: out<=0;
   37329: out<=1;
   37330: out<=0;
   37331: out<=1;
   37332: out<=1;
   37333: out<=1;
   37334: out<=0;
   37335: out<=0;
   37336: out<=1;
   37337: out<=1;
   37338: out<=1;
   37339: out<=1;
   37340: out<=0;
   37341: out<=1;
   37342: out<=1;
   37343: out<=0;
   37344: out<=0;
   37345: out<=1;
   37346: out<=1;
   37347: out<=0;
   37348: out<=1;
   37349: out<=1;
   37350: out<=1;
   37351: out<=1;
   37352: out<=0;
   37353: out<=0;
   37354: out<=1;
   37355: out<=1;
   37356: out<=1;
   37357: out<=0;
   37358: out<=1;
   37359: out<=0;
   37360: out<=0;
   37361: out<=0;
   37362: out<=0;
   37363: out<=0;
   37364: out<=0;
   37365: out<=1;
   37366: out<=1;
   37367: out<=0;
   37368: out<=1;
   37369: out<=0;
   37370: out<=1;
   37371: out<=0;
   37372: out<=1;
   37373: out<=1;
   37374: out<=0;
   37375: out<=0;
   37376: out<=0;
   37377: out<=0;
   37378: out<=0;
   37379: out<=0;
   37380: out<=0;
   37381: out<=1;
   37382: out<=1;
   37383: out<=0;
   37384: out<=1;
   37385: out<=0;
   37386: out<=1;
   37387: out<=0;
   37388: out<=1;
   37389: out<=1;
   37390: out<=0;
   37391: out<=0;
   37392: out<=0;
   37393: out<=1;
   37394: out<=1;
   37395: out<=0;
   37396: out<=1;
   37397: out<=1;
   37398: out<=1;
   37399: out<=1;
   37400: out<=0;
   37401: out<=0;
   37402: out<=1;
   37403: out<=1;
   37404: out<=1;
   37405: out<=0;
   37406: out<=1;
   37407: out<=0;
   37408: out<=0;
   37409: out<=1;
   37410: out<=0;
   37411: out<=1;
   37412: out<=1;
   37413: out<=1;
   37414: out<=0;
   37415: out<=0;
   37416: out<=1;
   37417: out<=1;
   37418: out<=1;
   37419: out<=1;
   37420: out<=0;
   37421: out<=1;
   37422: out<=1;
   37423: out<=0;
   37424: out<=0;
   37425: out<=0;
   37426: out<=1;
   37427: out<=1;
   37428: out<=0;
   37429: out<=1;
   37430: out<=0;
   37431: out<=1;
   37432: out<=0;
   37433: out<=1;
   37434: out<=1;
   37435: out<=0;
   37436: out<=0;
   37437: out<=0;
   37438: out<=0;
   37439: out<=0;
   37440: out<=1;
   37441: out<=1;
   37442: out<=1;
   37443: out<=1;
   37444: out<=1;
   37445: out<=0;
   37446: out<=0;
   37447: out<=1;
   37448: out<=0;
   37449: out<=1;
   37450: out<=0;
   37451: out<=1;
   37452: out<=0;
   37453: out<=0;
   37454: out<=1;
   37455: out<=1;
   37456: out<=0;
   37457: out<=1;
   37458: out<=1;
   37459: out<=0;
   37460: out<=1;
   37461: out<=1;
   37462: out<=1;
   37463: out<=1;
   37464: out<=0;
   37465: out<=0;
   37466: out<=1;
   37467: out<=1;
   37468: out<=1;
   37469: out<=0;
   37470: out<=1;
   37471: out<=0;
   37472: out<=0;
   37473: out<=1;
   37474: out<=0;
   37475: out<=1;
   37476: out<=1;
   37477: out<=1;
   37478: out<=0;
   37479: out<=0;
   37480: out<=1;
   37481: out<=1;
   37482: out<=1;
   37483: out<=1;
   37484: out<=0;
   37485: out<=1;
   37486: out<=1;
   37487: out<=0;
   37488: out<=1;
   37489: out<=1;
   37490: out<=0;
   37491: out<=0;
   37492: out<=1;
   37493: out<=0;
   37494: out<=1;
   37495: out<=0;
   37496: out<=1;
   37497: out<=0;
   37498: out<=0;
   37499: out<=1;
   37500: out<=1;
   37501: out<=1;
   37502: out<=1;
   37503: out<=1;
   37504: out<=0;
   37505: out<=0;
   37506: out<=0;
   37507: out<=0;
   37508: out<=0;
   37509: out<=1;
   37510: out<=1;
   37511: out<=0;
   37512: out<=1;
   37513: out<=0;
   37514: out<=1;
   37515: out<=0;
   37516: out<=1;
   37517: out<=1;
   37518: out<=0;
   37519: out<=0;
   37520: out<=1;
   37521: out<=0;
   37522: out<=0;
   37523: out<=1;
   37524: out<=0;
   37525: out<=0;
   37526: out<=0;
   37527: out<=0;
   37528: out<=1;
   37529: out<=1;
   37530: out<=0;
   37531: out<=0;
   37532: out<=0;
   37533: out<=1;
   37534: out<=0;
   37535: out<=1;
   37536: out<=0;
   37537: out<=1;
   37538: out<=0;
   37539: out<=1;
   37540: out<=1;
   37541: out<=1;
   37542: out<=0;
   37543: out<=0;
   37544: out<=1;
   37545: out<=1;
   37546: out<=1;
   37547: out<=1;
   37548: out<=0;
   37549: out<=1;
   37550: out<=1;
   37551: out<=0;
   37552: out<=1;
   37553: out<=1;
   37554: out<=0;
   37555: out<=0;
   37556: out<=1;
   37557: out<=0;
   37558: out<=1;
   37559: out<=0;
   37560: out<=1;
   37561: out<=0;
   37562: out<=0;
   37563: out<=1;
   37564: out<=1;
   37565: out<=1;
   37566: out<=1;
   37567: out<=1;
   37568: out<=1;
   37569: out<=1;
   37570: out<=1;
   37571: out<=1;
   37572: out<=1;
   37573: out<=0;
   37574: out<=0;
   37575: out<=1;
   37576: out<=0;
   37577: out<=1;
   37578: out<=0;
   37579: out<=1;
   37580: out<=0;
   37581: out<=0;
   37582: out<=1;
   37583: out<=1;
   37584: out<=1;
   37585: out<=0;
   37586: out<=0;
   37587: out<=1;
   37588: out<=0;
   37589: out<=0;
   37590: out<=0;
   37591: out<=0;
   37592: out<=1;
   37593: out<=1;
   37594: out<=0;
   37595: out<=0;
   37596: out<=0;
   37597: out<=1;
   37598: out<=0;
   37599: out<=1;
   37600: out<=0;
   37601: out<=1;
   37602: out<=0;
   37603: out<=1;
   37604: out<=1;
   37605: out<=1;
   37606: out<=0;
   37607: out<=0;
   37608: out<=1;
   37609: out<=1;
   37610: out<=1;
   37611: out<=1;
   37612: out<=0;
   37613: out<=1;
   37614: out<=1;
   37615: out<=0;
   37616: out<=0;
   37617: out<=0;
   37618: out<=1;
   37619: out<=1;
   37620: out<=0;
   37621: out<=1;
   37622: out<=0;
   37623: out<=1;
   37624: out<=0;
   37625: out<=1;
   37626: out<=1;
   37627: out<=0;
   37628: out<=0;
   37629: out<=0;
   37630: out<=0;
   37631: out<=0;
   37632: out<=0;
   37633: out<=1;
   37634: out<=1;
   37635: out<=0;
   37636: out<=1;
   37637: out<=1;
   37638: out<=1;
   37639: out<=1;
   37640: out<=0;
   37641: out<=0;
   37642: out<=1;
   37643: out<=1;
   37644: out<=1;
   37645: out<=0;
   37646: out<=1;
   37647: out<=0;
   37648: out<=1;
   37649: out<=1;
   37650: out<=1;
   37651: out<=1;
   37652: out<=1;
   37653: out<=0;
   37654: out<=0;
   37655: out<=1;
   37656: out<=0;
   37657: out<=1;
   37658: out<=0;
   37659: out<=1;
   37660: out<=0;
   37661: out<=0;
   37662: out<=1;
   37663: out<=1;
   37664: out<=1;
   37665: out<=1;
   37666: out<=0;
   37667: out<=0;
   37668: out<=1;
   37669: out<=0;
   37670: out<=1;
   37671: out<=0;
   37672: out<=1;
   37673: out<=0;
   37674: out<=0;
   37675: out<=1;
   37676: out<=1;
   37677: out<=1;
   37678: out<=1;
   37679: out<=1;
   37680: out<=0;
   37681: out<=1;
   37682: out<=0;
   37683: out<=1;
   37684: out<=1;
   37685: out<=1;
   37686: out<=0;
   37687: out<=0;
   37688: out<=1;
   37689: out<=1;
   37690: out<=1;
   37691: out<=1;
   37692: out<=0;
   37693: out<=1;
   37694: out<=1;
   37695: out<=0;
   37696: out<=0;
   37697: out<=1;
   37698: out<=1;
   37699: out<=0;
   37700: out<=1;
   37701: out<=1;
   37702: out<=1;
   37703: out<=1;
   37704: out<=0;
   37705: out<=0;
   37706: out<=1;
   37707: out<=1;
   37708: out<=1;
   37709: out<=0;
   37710: out<=1;
   37711: out<=0;
   37712: out<=0;
   37713: out<=0;
   37714: out<=0;
   37715: out<=0;
   37716: out<=0;
   37717: out<=1;
   37718: out<=1;
   37719: out<=0;
   37720: out<=1;
   37721: out<=0;
   37722: out<=1;
   37723: out<=0;
   37724: out<=1;
   37725: out<=1;
   37726: out<=0;
   37727: out<=0;
   37728: out<=0;
   37729: out<=0;
   37730: out<=1;
   37731: out<=1;
   37732: out<=0;
   37733: out<=1;
   37734: out<=0;
   37735: out<=1;
   37736: out<=0;
   37737: out<=1;
   37738: out<=1;
   37739: out<=0;
   37740: out<=0;
   37741: out<=0;
   37742: out<=0;
   37743: out<=0;
   37744: out<=0;
   37745: out<=1;
   37746: out<=0;
   37747: out<=1;
   37748: out<=1;
   37749: out<=1;
   37750: out<=0;
   37751: out<=0;
   37752: out<=1;
   37753: out<=1;
   37754: out<=1;
   37755: out<=1;
   37756: out<=0;
   37757: out<=1;
   37758: out<=1;
   37759: out<=0;
   37760: out<=1;
   37761: out<=0;
   37762: out<=0;
   37763: out<=1;
   37764: out<=0;
   37765: out<=0;
   37766: out<=0;
   37767: out<=0;
   37768: out<=1;
   37769: out<=1;
   37770: out<=0;
   37771: out<=0;
   37772: out<=0;
   37773: out<=1;
   37774: out<=0;
   37775: out<=1;
   37776: out<=1;
   37777: out<=1;
   37778: out<=1;
   37779: out<=1;
   37780: out<=1;
   37781: out<=0;
   37782: out<=0;
   37783: out<=1;
   37784: out<=0;
   37785: out<=1;
   37786: out<=0;
   37787: out<=1;
   37788: out<=0;
   37789: out<=0;
   37790: out<=1;
   37791: out<=1;
   37792: out<=0;
   37793: out<=0;
   37794: out<=1;
   37795: out<=1;
   37796: out<=0;
   37797: out<=1;
   37798: out<=0;
   37799: out<=1;
   37800: out<=0;
   37801: out<=1;
   37802: out<=1;
   37803: out<=0;
   37804: out<=0;
   37805: out<=0;
   37806: out<=0;
   37807: out<=0;
   37808: out<=0;
   37809: out<=1;
   37810: out<=0;
   37811: out<=1;
   37812: out<=1;
   37813: out<=1;
   37814: out<=0;
   37815: out<=0;
   37816: out<=1;
   37817: out<=1;
   37818: out<=1;
   37819: out<=1;
   37820: out<=0;
   37821: out<=1;
   37822: out<=1;
   37823: out<=0;
   37824: out<=1;
   37825: out<=0;
   37826: out<=0;
   37827: out<=1;
   37828: out<=0;
   37829: out<=0;
   37830: out<=0;
   37831: out<=0;
   37832: out<=1;
   37833: out<=1;
   37834: out<=0;
   37835: out<=0;
   37836: out<=0;
   37837: out<=1;
   37838: out<=0;
   37839: out<=1;
   37840: out<=0;
   37841: out<=0;
   37842: out<=0;
   37843: out<=0;
   37844: out<=0;
   37845: out<=1;
   37846: out<=1;
   37847: out<=0;
   37848: out<=1;
   37849: out<=0;
   37850: out<=1;
   37851: out<=0;
   37852: out<=1;
   37853: out<=1;
   37854: out<=0;
   37855: out<=0;
   37856: out<=1;
   37857: out<=1;
   37858: out<=0;
   37859: out<=0;
   37860: out<=1;
   37861: out<=0;
   37862: out<=1;
   37863: out<=0;
   37864: out<=1;
   37865: out<=0;
   37866: out<=0;
   37867: out<=1;
   37868: out<=1;
   37869: out<=1;
   37870: out<=1;
   37871: out<=1;
   37872: out<=0;
   37873: out<=1;
   37874: out<=0;
   37875: out<=1;
   37876: out<=1;
   37877: out<=1;
   37878: out<=0;
   37879: out<=0;
   37880: out<=1;
   37881: out<=1;
   37882: out<=1;
   37883: out<=1;
   37884: out<=0;
   37885: out<=1;
   37886: out<=1;
   37887: out<=0;
   37888: out<=0;
   37889: out<=0;
   37890: out<=1;
   37891: out<=1;
   37892: out<=1;
   37893: out<=0;
   37894: out<=1;
   37895: out<=0;
   37896: out<=1;
   37897: out<=0;
   37898: out<=0;
   37899: out<=1;
   37900: out<=0;
   37901: out<=0;
   37902: out<=0;
   37903: out<=0;
   37904: out<=1;
   37905: out<=0;
   37906: out<=1;
   37907: out<=0;
   37908: out<=1;
   37909: out<=1;
   37910: out<=0;
   37911: out<=0;
   37912: out<=1;
   37913: out<=1;
   37914: out<=1;
   37915: out<=1;
   37916: out<=1;
   37917: out<=0;
   37918: out<=0;
   37919: out<=1;
   37920: out<=0;
   37921: out<=1;
   37922: out<=1;
   37923: out<=0;
   37924: out<=0;
   37925: out<=0;
   37926: out<=0;
   37927: out<=0;
   37928: out<=1;
   37929: out<=1;
   37930: out<=0;
   37931: out<=0;
   37932: out<=1;
   37933: out<=0;
   37934: out<=1;
   37935: out<=0;
   37936: out<=1;
   37937: out<=1;
   37938: out<=1;
   37939: out<=1;
   37940: out<=0;
   37941: out<=1;
   37942: out<=1;
   37943: out<=0;
   37944: out<=1;
   37945: out<=0;
   37946: out<=1;
   37947: out<=0;
   37948: out<=0;
   37949: out<=0;
   37950: out<=1;
   37951: out<=1;
   37952: out<=1;
   37953: out<=1;
   37954: out<=0;
   37955: out<=0;
   37956: out<=0;
   37957: out<=1;
   37958: out<=0;
   37959: out<=1;
   37960: out<=0;
   37961: out<=1;
   37962: out<=1;
   37963: out<=0;
   37964: out<=1;
   37965: out<=1;
   37966: out<=1;
   37967: out<=1;
   37968: out<=1;
   37969: out<=0;
   37970: out<=1;
   37971: out<=0;
   37972: out<=1;
   37973: out<=1;
   37974: out<=0;
   37975: out<=0;
   37976: out<=1;
   37977: out<=1;
   37978: out<=1;
   37979: out<=1;
   37980: out<=1;
   37981: out<=0;
   37982: out<=0;
   37983: out<=1;
   37984: out<=0;
   37985: out<=1;
   37986: out<=1;
   37987: out<=0;
   37988: out<=0;
   37989: out<=0;
   37990: out<=0;
   37991: out<=0;
   37992: out<=1;
   37993: out<=1;
   37994: out<=0;
   37995: out<=0;
   37996: out<=1;
   37997: out<=0;
   37998: out<=1;
   37999: out<=0;
   38000: out<=0;
   38001: out<=0;
   38002: out<=0;
   38003: out<=0;
   38004: out<=1;
   38005: out<=0;
   38006: out<=0;
   38007: out<=1;
   38008: out<=0;
   38009: out<=1;
   38010: out<=0;
   38011: out<=1;
   38012: out<=1;
   38013: out<=1;
   38014: out<=0;
   38015: out<=0;
   38016: out<=1;
   38017: out<=1;
   38018: out<=0;
   38019: out<=0;
   38020: out<=0;
   38021: out<=1;
   38022: out<=0;
   38023: out<=1;
   38024: out<=0;
   38025: out<=1;
   38026: out<=1;
   38027: out<=0;
   38028: out<=1;
   38029: out<=1;
   38030: out<=1;
   38031: out<=1;
   38032: out<=1;
   38033: out<=0;
   38034: out<=1;
   38035: out<=0;
   38036: out<=1;
   38037: out<=1;
   38038: out<=0;
   38039: out<=0;
   38040: out<=1;
   38041: out<=1;
   38042: out<=1;
   38043: out<=1;
   38044: out<=1;
   38045: out<=0;
   38046: out<=0;
   38047: out<=1;
   38048: out<=1;
   38049: out<=0;
   38050: out<=0;
   38051: out<=1;
   38052: out<=1;
   38053: out<=1;
   38054: out<=1;
   38055: out<=1;
   38056: out<=0;
   38057: out<=0;
   38058: out<=1;
   38059: out<=1;
   38060: out<=0;
   38061: out<=1;
   38062: out<=0;
   38063: out<=1;
   38064: out<=1;
   38065: out<=1;
   38066: out<=1;
   38067: out<=1;
   38068: out<=0;
   38069: out<=1;
   38070: out<=1;
   38071: out<=0;
   38072: out<=1;
   38073: out<=0;
   38074: out<=1;
   38075: out<=0;
   38076: out<=0;
   38077: out<=0;
   38078: out<=1;
   38079: out<=1;
   38080: out<=0;
   38081: out<=0;
   38082: out<=1;
   38083: out<=1;
   38084: out<=1;
   38085: out<=0;
   38086: out<=1;
   38087: out<=0;
   38088: out<=1;
   38089: out<=0;
   38090: out<=0;
   38091: out<=1;
   38092: out<=0;
   38093: out<=0;
   38094: out<=0;
   38095: out<=0;
   38096: out<=1;
   38097: out<=0;
   38098: out<=1;
   38099: out<=0;
   38100: out<=1;
   38101: out<=1;
   38102: out<=0;
   38103: out<=0;
   38104: out<=1;
   38105: out<=1;
   38106: out<=1;
   38107: out<=1;
   38108: out<=1;
   38109: out<=0;
   38110: out<=0;
   38111: out<=1;
   38112: out<=1;
   38113: out<=0;
   38114: out<=0;
   38115: out<=1;
   38116: out<=1;
   38117: out<=1;
   38118: out<=1;
   38119: out<=1;
   38120: out<=0;
   38121: out<=0;
   38122: out<=1;
   38123: out<=1;
   38124: out<=0;
   38125: out<=1;
   38126: out<=0;
   38127: out<=1;
   38128: out<=0;
   38129: out<=0;
   38130: out<=0;
   38131: out<=0;
   38132: out<=1;
   38133: out<=0;
   38134: out<=0;
   38135: out<=1;
   38136: out<=0;
   38137: out<=1;
   38138: out<=0;
   38139: out<=1;
   38140: out<=1;
   38141: out<=1;
   38142: out<=0;
   38143: out<=0;
   38144: out<=1;
   38145: out<=0;
   38146: out<=1;
   38147: out<=0;
   38148: out<=1;
   38149: out<=1;
   38150: out<=0;
   38151: out<=0;
   38152: out<=1;
   38153: out<=1;
   38154: out<=1;
   38155: out<=1;
   38156: out<=1;
   38157: out<=0;
   38158: out<=0;
   38159: out<=1;
   38160: out<=1;
   38161: out<=1;
   38162: out<=0;
   38163: out<=0;
   38164: out<=0;
   38165: out<=1;
   38166: out<=0;
   38167: out<=1;
   38168: out<=0;
   38169: out<=1;
   38170: out<=1;
   38171: out<=0;
   38172: out<=1;
   38173: out<=1;
   38174: out<=1;
   38175: out<=1;
   38176: out<=0;
   38177: out<=0;
   38178: out<=0;
   38179: out<=0;
   38180: out<=1;
   38181: out<=0;
   38182: out<=0;
   38183: out<=1;
   38184: out<=0;
   38185: out<=1;
   38186: out<=0;
   38187: out<=1;
   38188: out<=1;
   38189: out<=1;
   38190: out<=0;
   38191: out<=0;
   38192: out<=0;
   38193: out<=1;
   38194: out<=1;
   38195: out<=0;
   38196: out<=0;
   38197: out<=0;
   38198: out<=0;
   38199: out<=0;
   38200: out<=1;
   38201: out<=1;
   38202: out<=0;
   38203: out<=0;
   38204: out<=1;
   38205: out<=0;
   38206: out<=1;
   38207: out<=0;
   38208: out<=1;
   38209: out<=0;
   38210: out<=1;
   38211: out<=0;
   38212: out<=1;
   38213: out<=1;
   38214: out<=0;
   38215: out<=0;
   38216: out<=1;
   38217: out<=1;
   38218: out<=1;
   38219: out<=1;
   38220: out<=1;
   38221: out<=0;
   38222: out<=0;
   38223: out<=1;
   38224: out<=0;
   38225: out<=0;
   38226: out<=1;
   38227: out<=1;
   38228: out<=1;
   38229: out<=0;
   38230: out<=1;
   38231: out<=0;
   38232: out<=1;
   38233: out<=0;
   38234: out<=0;
   38235: out<=1;
   38236: out<=0;
   38237: out<=0;
   38238: out<=0;
   38239: out<=0;
   38240: out<=1;
   38241: out<=1;
   38242: out<=1;
   38243: out<=1;
   38244: out<=0;
   38245: out<=1;
   38246: out<=1;
   38247: out<=0;
   38248: out<=1;
   38249: out<=0;
   38250: out<=1;
   38251: out<=0;
   38252: out<=0;
   38253: out<=0;
   38254: out<=1;
   38255: out<=1;
   38256: out<=0;
   38257: out<=1;
   38258: out<=1;
   38259: out<=0;
   38260: out<=0;
   38261: out<=0;
   38262: out<=0;
   38263: out<=0;
   38264: out<=1;
   38265: out<=1;
   38266: out<=0;
   38267: out<=0;
   38268: out<=1;
   38269: out<=0;
   38270: out<=1;
   38271: out<=0;
   38272: out<=1;
   38273: out<=0;
   38274: out<=1;
   38275: out<=0;
   38276: out<=1;
   38277: out<=1;
   38278: out<=0;
   38279: out<=0;
   38280: out<=1;
   38281: out<=1;
   38282: out<=1;
   38283: out<=1;
   38284: out<=1;
   38285: out<=0;
   38286: out<=0;
   38287: out<=1;
   38288: out<=0;
   38289: out<=0;
   38290: out<=1;
   38291: out<=1;
   38292: out<=1;
   38293: out<=0;
   38294: out<=1;
   38295: out<=0;
   38296: out<=1;
   38297: out<=0;
   38298: out<=0;
   38299: out<=1;
   38300: out<=0;
   38301: out<=0;
   38302: out<=0;
   38303: out<=0;
   38304: out<=0;
   38305: out<=0;
   38306: out<=0;
   38307: out<=0;
   38308: out<=1;
   38309: out<=0;
   38310: out<=0;
   38311: out<=1;
   38312: out<=0;
   38313: out<=1;
   38314: out<=0;
   38315: out<=1;
   38316: out<=1;
   38317: out<=1;
   38318: out<=0;
   38319: out<=0;
   38320: out<=1;
   38321: out<=0;
   38322: out<=0;
   38323: out<=1;
   38324: out<=1;
   38325: out<=1;
   38326: out<=1;
   38327: out<=1;
   38328: out<=0;
   38329: out<=0;
   38330: out<=1;
   38331: out<=1;
   38332: out<=0;
   38333: out<=1;
   38334: out<=0;
   38335: out<=1;
   38336: out<=1;
   38337: out<=0;
   38338: out<=1;
   38339: out<=0;
   38340: out<=1;
   38341: out<=1;
   38342: out<=0;
   38343: out<=0;
   38344: out<=1;
   38345: out<=1;
   38346: out<=1;
   38347: out<=1;
   38348: out<=1;
   38349: out<=0;
   38350: out<=0;
   38351: out<=1;
   38352: out<=1;
   38353: out<=1;
   38354: out<=0;
   38355: out<=0;
   38356: out<=0;
   38357: out<=1;
   38358: out<=0;
   38359: out<=1;
   38360: out<=0;
   38361: out<=1;
   38362: out<=1;
   38363: out<=0;
   38364: out<=1;
   38365: out<=1;
   38366: out<=1;
   38367: out<=1;
   38368: out<=1;
   38369: out<=1;
   38370: out<=1;
   38371: out<=1;
   38372: out<=0;
   38373: out<=1;
   38374: out<=1;
   38375: out<=0;
   38376: out<=1;
   38377: out<=0;
   38378: out<=1;
   38379: out<=0;
   38380: out<=0;
   38381: out<=0;
   38382: out<=1;
   38383: out<=1;
   38384: out<=1;
   38385: out<=0;
   38386: out<=0;
   38387: out<=1;
   38388: out<=1;
   38389: out<=1;
   38390: out<=1;
   38391: out<=1;
   38392: out<=0;
   38393: out<=0;
   38394: out<=1;
   38395: out<=1;
   38396: out<=0;
   38397: out<=1;
   38398: out<=0;
   38399: out<=1;
   38400: out<=1;
   38401: out<=0;
   38402: out<=0;
   38403: out<=1;
   38404: out<=1;
   38405: out<=1;
   38406: out<=1;
   38407: out<=1;
   38408: out<=0;
   38409: out<=0;
   38410: out<=1;
   38411: out<=1;
   38412: out<=0;
   38413: out<=1;
   38414: out<=0;
   38415: out<=1;
   38416: out<=1;
   38417: out<=1;
   38418: out<=1;
   38419: out<=1;
   38420: out<=0;
   38421: out<=1;
   38422: out<=1;
   38423: out<=0;
   38424: out<=1;
   38425: out<=0;
   38426: out<=1;
   38427: out<=0;
   38428: out<=0;
   38429: out<=0;
   38430: out<=1;
   38431: out<=1;
   38432: out<=1;
   38433: out<=1;
   38434: out<=0;
   38435: out<=0;
   38436: out<=0;
   38437: out<=1;
   38438: out<=0;
   38439: out<=1;
   38440: out<=0;
   38441: out<=1;
   38442: out<=1;
   38443: out<=0;
   38444: out<=1;
   38445: out<=1;
   38446: out<=1;
   38447: out<=1;
   38448: out<=1;
   38449: out<=0;
   38450: out<=1;
   38451: out<=0;
   38452: out<=1;
   38453: out<=1;
   38454: out<=0;
   38455: out<=0;
   38456: out<=1;
   38457: out<=1;
   38458: out<=1;
   38459: out<=1;
   38460: out<=1;
   38461: out<=0;
   38462: out<=0;
   38463: out<=1;
   38464: out<=1;
   38465: out<=0;
   38466: out<=0;
   38467: out<=1;
   38468: out<=1;
   38469: out<=1;
   38470: out<=1;
   38471: out<=1;
   38472: out<=0;
   38473: out<=0;
   38474: out<=1;
   38475: out<=1;
   38476: out<=0;
   38477: out<=1;
   38478: out<=0;
   38479: out<=1;
   38480: out<=0;
   38481: out<=0;
   38482: out<=0;
   38483: out<=0;
   38484: out<=1;
   38485: out<=0;
   38486: out<=0;
   38487: out<=1;
   38488: out<=0;
   38489: out<=1;
   38490: out<=0;
   38491: out<=1;
   38492: out<=1;
   38493: out<=1;
   38494: out<=0;
   38495: out<=0;
   38496: out<=0;
   38497: out<=0;
   38498: out<=1;
   38499: out<=1;
   38500: out<=1;
   38501: out<=0;
   38502: out<=1;
   38503: out<=0;
   38504: out<=1;
   38505: out<=0;
   38506: out<=0;
   38507: out<=1;
   38508: out<=0;
   38509: out<=0;
   38510: out<=0;
   38511: out<=0;
   38512: out<=1;
   38513: out<=0;
   38514: out<=1;
   38515: out<=0;
   38516: out<=1;
   38517: out<=1;
   38518: out<=0;
   38519: out<=0;
   38520: out<=1;
   38521: out<=1;
   38522: out<=1;
   38523: out<=1;
   38524: out<=1;
   38525: out<=0;
   38526: out<=0;
   38527: out<=1;
   38528: out<=0;
   38529: out<=1;
   38530: out<=1;
   38531: out<=0;
   38532: out<=0;
   38533: out<=0;
   38534: out<=0;
   38535: out<=0;
   38536: out<=1;
   38537: out<=1;
   38538: out<=0;
   38539: out<=0;
   38540: out<=1;
   38541: out<=0;
   38542: out<=1;
   38543: out<=0;
   38544: out<=1;
   38545: out<=1;
   38546: out<=1;
   38547: out<=1;
   38548: out<=0;
   38549: out<=1;
   38550: out<=1;
   38551: out<=0;
   38552: out<=1;
   38553: out<=0;
   38554: out<=1;
   38555: out<=0;
   38556: out<=0;
   38557: out<=0;
   38558: out<=1;
   38559: out<=1;
   38560: out<=0;
   38561: out<=0;
   38562: out<=1;
   38563: out<=1;
   38564: out<=1;
   38565: out<=0;
   38566: out<=1;
   38567: out<=0;
   38568: out<=1;
   38569: out<=0;
   38570: out<=0;
   38571: out<=1;
   38572: out<=0;
   38573: out<=0;
   38574: out<=0;
   38575: out<=0;
   38576: out<=1;
   38577: out<=0;
   38578: out<=1;
   38579: out<=0;
   38580: out<=1;
   38581: out<=1;
   38582: out<=0;
   38583: out<=0;
   38584: out<=1;
   38585: out<=1;
   38586: out<=1;
   38587: out<=1;
   38588: out<=1;
   38589: out<=0;
   38590: out<=0;
   38591: out<=1;
   38592: out<=0;
   38593: out<=1;
   38594: out<=1;
   38595: out<=0;
   38596: out<=0;
   38597: out<=0;
   38598: out<=0;
   38599: out<=0;
   38600: out<=1;
   38601: out<=1;
   38602: out<=0;
   38603: out<=0;
   38604: out<=1;
   38605: out<=0;
   38606: out<=1;
   38607: out<=0;
   38608: out<=0;
   38609: out<=0;
   38610: out<=0;
   38611: out<=0;
   38612: out<=1;
   38613: out<=0;
   38614: out<=0;
   38615: out<=1;
   38616: out<=0;
   38617: out<=1;
   38618: out<=0;
   38619: out<=1;
   38620: out<=1;
   38621: out<=1;
   38622: out<=0;
   38623: out<=0;
   38624: out<=1;
   38625: out<=1;
   38626: out<=0;
   38627: out<=0;
   38628: out<=0;
   38629: out<=1;
   38630: out<=0;
   38631: out<=1;
   38632: out<=0;
   38633: out<=1;
   38634: out<=1;
   38635: out<=0;
   38636: out<=1;
   38637: out<=1;
   38638: out<=1;
   38639: out<=1;
   38640: out<=1;
   38641: out<=0;
   38642: out<=1;
   38643: out<=0;
   38644: out<=1;
   38645: out<=1;
   38646: out<=0;
   38647: out<=0;
   38648: out<=1;
   38649: out<=1;
   38650: out<=1;
   38651: out<=1;
   38652: out<=1;
   38653: out<=0;
   38654: out<=0;
   38655: out<=1;
   38656: out<=0;
   38657: out<=0;
   38658: out<=0;
   38659: out<=0;
   38660: out<=1;
   38661: out<=0;
   38662: out<=0;
   38663: out<=1;
   38664: out<=0;
   38665: out<=1;
   38666: out<=0;
   38667: out<=1;
   38668: out<=1;
   38669: out<=1;
   38670: out<=0;
   38671: out<=0;
   38672: out<=1;
   38673: out<=0;
   38674: out<=0;
   38675: out<=1;
   38676: out<=1;
   38677: out<=1;
   38678: out<=1;
   38679: out<=1;
   38680: out<=0;
   38681: out<=0;
   38682: out<=1;
   38683: out<=1;
   38684: out<=0;
   38685: out<=1;
   38686: out<=0;
   38687: out<=1;
   38688: out<=1;
   38689: out<=0;
   38690: out<=1;
   38691: out<=0;
   38692: out<=1;
   38693: out<=1;
   38694: out<=0;
   38695: out<=0;
   38696: out<=1;
   38697: out<=1;
   38698: out<=1;
   38699: out<=1;
   38700: out<=1;
   38701: out<=0;
   38702: out<=0;
   38703: out<=1;
   38704: out<=0;
   38705: out<=0;
   38706: out<=1;
   38707: out<=1;
   38708: out<=1;
   38709: out<=0;
   38710: out<=1;
   38711: out<=0;
   38712: out<=1;
   38713: out<=0;
   38714: out<=0;
   38715: out<=1;
   38716: out<=0;
   38717: out<=0;
   38718: out<=0;
   38719: out<=0;
   38720: out<=1;
   38721: out<=1;
   38722: out<=1;
   38723: out<=1;
   38724: out<=0;
   38725: out<=1;
   38726: out<=1;
   38727: out<=0;
   38728: out<=1;
   38729: out<=0;
   38730: out<=1;
   38731: out<=0;
   38732: out<=0;
   38733: out<=0;
   38734: out<=1;
   38735: out<=1;
   38736: out<=1;
   38737: out<=0;
   38738: out<=0;
   38739: out<=1;
   38740: out<=1;
   38741: out<=1;
   38742: out<=1;
   38743: out<=1;
   38744: out<=0;
   38745: out<=0;
   38746: out<=1;
   38747: out<=1;
   38748: out<=0;
   38749: out<=1;
   38750: out<=0;
   38751: out<=1;
   38752: out<=1;
   38753: out<=0;
   38754: out<=1;
   38755: out<=0;
   38756: out<=1;
   38757: out<=1;
   38758: out<=0;
   38759: out<=0;
   38760: out<=1;
   38761: out<=1;
   38762: out<=1;
   38763: out<=1;
   38764: out<=1;
   38765: out<=0;
   38766: out<=0;
   38767: out<=1;
   38768: out<=1;
   38769: out<=1;
   38770: out<=0;
   38771: out<=0;
   38772: out<=0;
   38773: out<=1;
   38774: out<=0;
   38775: out<=1;
   38776: out<=0;
   38777: out<=1;
   38778: out<=1;
   38779: out<=0;
   38780: out<=1;
   38781: out<=1;
   38782: out<=1;
   38783: out<=1;
   38784: out<=0;
   38785: out<=0;
   38786: out<=0;
   38787: out<=0;
   38788: out<=1;
   38789: out<=0;
   38790: out<=0;
   38791: out<=1;
   38792: out<=0;
   38793: out<=1;
   38794: out<=0;
   38795: out<=1;
   38796: out<=1;
   38797: out<=1;
   38798: out<=0;
   38799: out<=0;
   38800: out<=0;
   38801: out<=1;
   38802: out<=1;
   38803: out<=0;
   38804: out<=0;
   38805: out<=0;
   38806: out<=0;
   38807: out<=0;
   38808: out<=1;
   38809: out<=1;
   38810: out<=0;
   38811: out<=0;
   38812: out<=1;
   38813: out<=0;
   38814: out<=1;
   38815: out<=0;
   38816: out<=1;
   38817: out<=0;
   38818: out<=1;
   38819: out<=0;
   38820: out<=1;
   38821: out<=1;
   38822: out<=0;
   38823: out<=0;
   38824: out<=1;
   38825: out<=1;
   38826: out<=1;
   38827: out<=1;
   38828: out<=1;
   38829: out<=0;
   38830: out<=0;
   38831: out<=1;
   38832: out<=1;
   38833: out<=1;
   38834: out<=0;
   38835: out<=0;
   38836: out<=0;
   38837: out<=1;
   38838: out<=0;
   38839: out<=1;
   38840: out<=0;
   38841: out<=1;
   38842: out<=1;
   38843: out<=0;
   38844: out<=1;
   38845: out<=1;
   38846: out<=1;
   38847: out<=1;
   38848: out<=1;
   38849: out<=1;
   38850: out<=1;
   38851: out<=1;
   38852: out<=0;
   38853: out<=1;
   38854: out<=1;
   38855: out<=0;
   38856: out<=1;
   38857: out<=0;
   38858: out<=1;
   38859: out<=0;
   38860: out<=0;
   38861: out<=0;
   38862: out<=1;
   38863: out<=1;
   38864: out<=0;
   38865: out<=1;
   38866: out<=1;
   38867: out<=0;
   38868: out<=0;
   38869: out<=0;
   38870: out<=0;
   38871: out<=0;
   38872: out<=1;
   38873: out<=1;
   38874: out<=0;
   38875: out<=0;
   38876: out<=1;
   38877: out<=0;
   38878: out<=1;
   38879: out<=0;
   38880: out<=1;
   38881: out<=0;
   38882: out<=1;
   38883: out<=0;
   38884: out<=1;
   38885: out<=1;
   38886: out<=0;
   38887: out<=0;
   38888: out<=1;
   38889: out<=1;
   38890: out<=1;
   38891: out<=1;
   38892: out<=1;
   38893: out<=0;
   38894: out<=0;
   38895: out<=1;
   38896: out<=0;
   38897: out<=0;
   38898: out<=1;
   38899: out<=1;
   38900: out<=1;
   38901: out<=0;
   38902: out<=1;
   38903: out<=0;
   38904: out<=1;
   38905: out<=0;
   38906: out<=0;
   38907: out<=1;
   38908: out<=0;
   38909: out<=0;
   38910: out<=0;
   38911: out<=0;
   38912: out<=0;
   38913: out<=0;
   38914: out<=0;
   38915: out<=0;
   38916: out<=1;
   38917: out<=0;
   38918: out<=0;
   38919: out<=1;
   38920: out<=1;
   38921: out<=0;
   38922: out<=1;
   38923: out<=0;
   38924: out<=0;
   38925: out<=0;
   38926: out<=1;
   38927: out<=1;
   38928: out<=1;
   38929: out<=0;
   38930: out<=0;
   38931: out<=1;
   38932: out<=1;
   38933: out<=1;
   38934: out<=1;
   38935: out<=1;
   38936: out<=1;
   38937: out<=1;
   38938: out<=0;
   38939: out<=0;
   38940: out<=1;
   38941: out<=0;
   38942: out<=1;
   38943: out<=0;
   38944: out<=0;
   38945: out<=1;
   38946: out<=0;
   38947: out<=1;
   38948: out<=0;
   38949: out<=0;
   38950: out<=1;
   38951: out<=1;
   38952: out<=1;
   38953: out<=1;
   38954: out<=1;
   38955: out<=1;
   38956: out<=1;
   38957: out<=0;
   38958: out<=0;
   38959: out<=1;
   38960: out<=1;
   38961: out<=1;
   38962: out<=0;
   38963: out<=0;
   38964: out<=0;
   38965: out<=1;
   38966: out<=0;
   38967: out<=1;
   38968: out<=1;
   38969: out<=0;
   38970: out<=0;
   38971: out<=1;
   38972: out<=0;
   38973: out<=0;
   38974: out<=0;
   38975: out<=0;
   38976: out<=1;
   38977: out<=1;
   38978: out<=1;
   38979: out<=1;
   38980: out<=0;
   38981: out<=1;
   38982: out<=1;
   38983: out<=0;
   38984: out<=0;
   38985: out<=1;
   38986: out<=0;
   38987: out<=1;
   38988: out<=1;
   38989: out<=1;
   38990: out<=0;
   38991: out<=0;
   38992: out<=1;
   38993: out<=0;
   38994: out<=0;
   38995: out<=1;
   38996: out<=1;
   38997: out<=1;
   38998: out<=1;
   38999: out<=1;
   39000: out<=1;
   39001: out<=1;
   39002: out<=0;
   39003: out<=0;
   39004: out<=1;
   39005: out<=0;
   39006: out<=1;
   39007: out<=0;
   39008: out<=0;
   39009: out<=1;
   39010: out<=0;
   39011: out<=1;
   39012: out<=0;
   39013: out<=0;
   39014: out<=1;
   39015: out<=1;
   39016: out<=1;
   39017: out<=1;
   39018: out<=1;
   39019: out<=1;
   39020: out<=1;
   39021: out<=0;
   39022: out<=0;
   39023: out<=1;
   39024: out<=0;
   39025: out<=0;
   39026: out<=1;
   39027: out<=1;
   39028: out<=1;
   39029: out<=0;
   39030: out<=1;
   39031: out<=0;
   39032: out<=0;
   39033: out<=1;
   39034: out<=1;
   39035: out<=0;
   39036: out<=1;
   39037: out<=1;
   39038: out<=1;
   39039: out<=1;
   39040: out<=0;
   39041: out<=0;
   39042: out<=0;
   39043: out<=0;
   39044: out<=1;
   39045: out<=0;
   39046: out<=0;
   39047: out<=1;
   39048: out<=1;
   39049: out<=0;
   39050: out<=1;
   39051: out<=0;
   39052: out<=0;
   39053: out<=0;
   39054: out<=1;
   39055: out<=1;
   39056: out<=0;
   39057: out<=1;
   39058: out<=1;
   39059: out<=0;
   39060: out<=0;
   39061: out<=0;
   39062: out<=0;
   39063: out<=0;
   39064: out<=0;
   39065: out<=0;
   39066: out<=1;
   39067: out<=1;
   39068: out<=0;
   39069: out<=1;
   39070: out<=0;
   39071: out<=1;
   39072: out<=0;
   39073: out<=1;
   39074: out<=0;
   39075: out<=1;
   39076: out<=0;
   39077: out<=0;
   39078: out<=1;
   39079: out<=1;
   39080: out<=1;
   39081: out<=1;
   39082: out<=1;
   39083: out<=1;
   39084: out<=1;
   39085: out<=0;
   39086: out<=0;
   39087: out<=1;
   39088: out<=0;
   39089: out<=0;
   39090: out<=1;
   39091: out<=1;
   39092: out<=1;
   39093: out<=0;
   39094: out<=1;
   39095: out<=0;
   39096: out<=0;
   39097: out<=1;
   39098: out<=1;
   39099: out<=0;
   39100: out<=1;
   39101: out<=1;
   39102: out<=1;
   39103: out<=1;
   39104: out<=1;
   39105: out<=1;
   39106: out<=1;
   39107: out<=1;
   39108: out<=0;
   39109: out<=1;
   39110: out<=1;
   39111: out<=0;
   39112: out<=0;
   39113: out<=1;
   39114: out<=0;
   39115: out<=1;
   39116: out<=1;
   39117: out<=1;
   39118: out<=0;
   39119: out<=0;
   39120: out<=0;
   39121: out<=1;
   39122: out<=1;
   39123: out<=0;
   39124: out<=0;
   39125: out<=0;
   39126: out<=0;
   39127: out<=0;
   39128: out<=0;
   39129: out<=0;
   39130: out<=1;
   39131: out<=1;
   39132: out<=0;
   39133: out<=1;
   39134: out<=0;
   39135: out<=1;
   39136: out<=0;
   39137: out<=1;
   39138: out<=0;
   39139: out<=1;
   39140: out<=0;
   39141: out<=0;
   39142: out<=1;
   39143: out<=1;
   39144: out<=1;
   39145: out<=1;
   39146: out<=1;
   39147: out<=1;
   39148: out<=1;
   39149: out<=0;
   39150: out<=0;
   39151: out<=1;
   39152: out<=1;
   39153: out<=1;
   39154: out<=0;
   39155: out<=0;
   39156: out<=0;
   39157: out<=1;
   39158: out<=0;
   39159: out<=1;
   39160: out<=1;
   39161: out<=0;
   39162: out<=0;
   39163: out<=1;
   39164: out<=0;
   39165: out<=0;
   39166: out<=0;
   39167: out<=0;
   39168: out<=1;
   39169: out<=0;
   39170: out<=0;
   39171: out<=1;
   39172: out<=1;
   39173: out<=1;
   39174: out<=1;
   39175: out<=1;
   39176: out<=1;
   39177: out<=1;
   39178: out<=0;
   39179: out<=0;
   39180: out<=1;
   39181: out<=0;
   39182: out<=1;
   39183: out<=0;
   39184: out<=1;
   39185: out<=1;
   39186: out<=1;
   39187: out<=1;
   39188: out<=0;
   39189: out<=1;
   39190: out<=1;
   39191: out<=0;
   39192: out<=0;
   39193: out<=1;
   39194: out<=0;
   39195: out<=1;
   39196: out<=1;
   39197: out<=1;
   39198: out<=0;
   39199: out<=0;
   39200: out<=0;
   39201: out<=0;
   39202: out<=1;
   39203: out<=1;
   39204: out<=1;
   39205: out<=0;
   39206: out<=1;
   39207: out<=0;
   39208: out<=0;
   39209: out<=1;
   39210: out<=1;
   39211: out<=0;
   39212: out<=1;
   39213: out<=1;
   39214: out<=1;
   39215: out<=1;
   39216: out<=0;
   39217: out<=1;
   39218: out<=0;
   39219: out<=1;
   39220: out<=0;
   39221: out<=0;
   39222: out<=1;
   39223: out<=1;
   39224: out<=1;
   39225: out<=1;
   39226: out<=1;
   39227: out<=1;
   39228: out<=1;
   39229: out<=0;
   39230: out<=0;
   39231: out<=1;
   39232: out<=1;
   39233: out<=0;
   39234: out<=0;
   39235: out<=1;
   39236: out<=1;
   39237: out<=1;
   39238: out<=1;
   39239: out<=1;
   39240: out<=1;
   39241: out<=1;
   39242: out<=0;
   39243: out<=0;
   39244: out<=1;
   39245: out<=0;
   39246: out<=1;
   39247: out<=0;
   39248: out<=0;
   39249: out<=0;
   39250: out<=0;
   39251: out<=0;
   39252: out<=1;
   39253: out<=0;
   39254: out<=0;
   39255: out<=1;
   39256: out<=1;
   39257: out<=0;
   39258: out<=1;
   39259: out<=0;
   39260: out<=0;
   39261: out<=0;
   39262: out<=1;
   39263: out<=1;
   39264: out<=1;
   39265: out<=1;
   39266: out<=0;
   39267: out<=0;
   39268: out<=0;
   39269: out<=1;
   39270: out<=0;
   39271: out<=1;
   39272: out<=1;
   39273: out<=0;
   39274: out<=0;
   39275: out<=1;
   39276: out<=0;
   39277: out<=0;
   39278: out<=0;
   39279: out<=0;
   39280: out<=0;
   39281: out<=1;
   39282: out<=0;
   39283: out<=1;
   39284: out<=0;
   39285: out<=0;
   39286: out<=1;
   39287: out<=1;
   39288: out<=1;
   39289: out<=1;
   39290: out<=1;
   39291: out<=1;
   39292: out<=1;
   39293: out<=0;
   39294: out<=0;
   39295: out<=1;
   39296: out<=0;
   39297: out<=1;
   39298: out<=1;
   39299: out<=0;
   39300: out<=0;
   39301: out<=0;
   39302: out<=0;
   39303: out<=0;
   39304: out<=0;
   39305: out<=0;
   39306: out<=1;
   39307: out<=1;
   39308: out<=0;
   39309: out<=1;
   39310: out<=0;
   39311: out<=1;
   39312: out<=1;
   39313: out<=1;
   39314: out<=1;
   39315: out<=1;
   39316: out<=0;
   39317: out<=1;
   39318: out<=1;
   39319: out<=0;
   39320: out<=0;
   39321: out<=1;
   39322: out<=0;
   39323: out<=1;
   39324: out<=1;
   39325: out<=1;
   39326: out<=0;
   39327: out<=0;
   39328: out<=1;
   39329: out<=1;
   39330: out<=0;
   39331: out<=0;
   39332: out<=0;
   39333: out<=1;
   39334: out<=0;
   39335: out<=1;
   39336: out<=1;
   39337: out<=0;
   39338: out<=0;
   39339: out<=1;
   39340: out<=0;
   39341: out<=0;
   39342: out<=0;
   39343: out<=0;
   39344: out<=0;
   39345: out<=1;
   39346: out<=0;
   39347: out<=1;
   39348: out<=0;
   39349: out<=0;
   39350: out<=1;
   39351: out<=1;
   39352: out<=1;
   39353: out<=1;
   39354: out<=1;
   39355: out<=1;
   39356: out<=1;
   39357: out<=0;
   39358: out<=0;
   39359: out<=1;
   39360: out<=0;
   39361: out<=1;
   39362: out<=1;
   39363: out<=0;
   39364: out<=0;
   39365: out<=0;
   39366: out<=0;
   39367: out<=0;
   39368: out<=0;
   39369: out<=0;
   39370: out<=1;
   39371: out<=1;
   39372: out<=0;
   39373: out<=1;
   39374: out<=0;
   39375: out<=1;
   39376: out<=0;
   39377: out<=0;
   39378: out<=0;
   39379: out<=0;
   39380: out<=1;
   39381: out<=0;
   39382: out<=0;
   39383: out<=1;
   39384: out<=1;
   39385: out<=0;
   39386: out<=1;
   39387: out<=0;
   39388: out<=0;
   39389: out<=0;
   39390: out<=1;
   39391: out<=1;
   39392: out<=0;
   39393: out<=0;
   39394: out<=1;
   39395: out<=1;
   39396: out<=1;
   39397: out<=0;
   39398: out<=1;
   39399: out<=0;
   39400: out<=0;
   39401: out<=1;
   39402: out<=1;
   39403: out<=0;
   39404: out<=1;
   39405: out<=1;
   39406: out<=1;
   39407: out<=1;
   39408: out<=0;
   39409: out<=1;
   39410: out<=0;
   39411: out<=1;
   39412: out<=0;
   39413: out<=0;
   39414: out<=1;
   39415: out<=1;
   39416: out<=1;
   39417: out<=1;
   39418: out<=1;
   39419: out<=1;
   39420: out<=1;
   39421: out<=0;
   39422: out<=0;
   39423: out<=1;
   39424: out<=0;
   39425: out<=1;
   39426: out<=0;
   39427: out<=1;
   39428: out<=0;
   39429: out<=0;
   39430: out<=1;
   39431: out<=1;
   39432: out<=1;
   39433: out<=1;
   39434: out<=1;
   39435: out<=1;
   39436: out<=1;
   39437: out<=0;
   39438: out<=0;
   39439: out<=1;
   39440: out<=0;
   39441: out<=0;
   39442: out<=1;
   39443: out<=1;
   39444: out<=1;
   39445: out<=0;
   39446: out<=1;
   39447: out<=0;
   39448: out<=0;
   39449: out<=1;
   39450: out<=1;
   39451: out<=0;
   39452: out<=1;
   39453: out<=1;
   39454: out<=1;
   39455: out<=1;
   39456: out<=0;
   39457: out<=0;
   39458: out<=0;
   39459: out<=0;
   39460: out<=1;
   39461: out<=0;
   39462: out<=0;
   39463: out<=1;
   39464: out<=1;
   39465: out<=0;
   39466: out<=1;
   39467: out<=0;
   39468: out<=0;
   39469: out<=0;
   39470: out<=1;
   39471: out<=1;
   39472: out<=0;
   39473: out<=1;
   39474: out<=1;
   39475: out<=0;
   39476: out<=0;
   39477: out<=0;
   39478: out<=0;
   39479: out<=0;
   39480: out<=0;
   39481: out<=0;
   39482: out<=1;
   39483: out<=1;
   39484: out<=0;
   39485: out<=1;
   39486: out<=0;
   39487: out<=1;
   39488: out<=0;
   39489: out<=1;
   39490: out<=0;
   39491: out<=1;
   39492: out<=0;
   39493: out<=0;
   39494: out<=1;
   39495: out<=1;
   39496: out<=1;
   39497: out<=1;
   39498: out<=1;
   39499: out<=1;
   39500: out<=1;
   39501: out<=0;
   39502: out<=0;
   39503: out<=1;
   39504: out<=1;
   39505: out<=1;
   39506: out<=0;
   39507: out<=0;
   39508: out<=0;
   39509: out<=1;
   39510: out<=0;
   39511: out<=1;
   39512: out<=1;
   39513: out<=0;
   39514: out<=0;
   39515: out<=1;
   39516: out<=0;
   39517: out<=0;
   39518: out<=0;
   39519: out<=0;
   39520: out<=1;
   39521: out<=1;
   39522: out<=1;
   39523: out<=1;
   39524: out<=0;
   39525: out<=1;
   39526: out<=1;
   39527: out<=0;
   39528: out<=0;
   39529: out<=1;
   39530: out<=0;
   39531: out<=1;
   39532: out<=1;
   39533: out<=1;
   39534: out<=0;
   39535: out<=0;
   39536: out<=0;
   39537: out<=1;
   39538: out<=1;
   39539: out<=0;
   39540: out<=0;
   39541: out<=0;
   39542: out<=0;
   39543: out<=0;
   39544: out<=0;
   39545: out<=0;
   39546: out<=1;
   39547: out<=1;
   39548: out<=0;
   39549: out<=1;
   39550: out<=0;
   39551: out<=1;
   39552: out<=0;
   39553: out<=1;
   39554: out<=0;
   39555: out<=1;
   39556: out<=0;
   39557: out<=0;
   39558: out<=1;
   39559: out<=1;
   39560: out<=1;
   39561: out<=1;
   39562: out<=1;
   39563: out<=1;
   39564: out<=1;
   39565: out<=0;
   39566: out<=0;
   39567: out<=1;
   39568: out<=1;
   39569: out<=1;
   39570: out<=0;
   39571: out<=0;
   39572: out<=0;
   39573: out<=1;
   39574: out<=0;
   39575: out<=1;
   39576: out<=1;
   39577: out<=0;
   39578: out<=0;
   39579: out<=1;
   39580: out<=0;
   39581: out<=0;
   39582: out<=0;
   39583: out<=0;
   39584: out<=0;
   39585: out<=0;
   39586: out<=0;
   39587: out<=0;
   39588: out<=1;
   39589: out<=0;
   39590: out<=0;
   39591: out<=1;
   39592: out<=1;
   39593: out<=0;
   39594: out<=1;
   39595: out<=0;
   39596: out<=0;
   39597: out<=0;
   39598: out<=1;
   39599: out<=1;
   39600: out<=1;
   39601: out<=0;
   39602: out<=0;
   39603: out<=1;
   39604: out<=1;
   39605: out<=1;
   39606: out<=1;
   39607: out<=1;
   39608: out<=1;
   39609: out<=1;
   39610: out<=0;
   39611: out<=0;
   39612: out<=1;
   39613: out<=0;
   39614: out<=1;
   39615: out<=0;
   39616: out<=0;
   39617: out<=1;
   39618: out<=0;
   39619: out<=1;
   39620: out<=0;
   39621: out<=0;
   39622: out<=1;
   39623: out<=1;
   39624: out<=1;
   39625: out<=1;
   39626: out<=1;
   39627: out<=1;
   39628: out<=1;
   39629: out<=0;
   39630: out<=0;
   39631: out<=1;
   39632: out<=0;
   39633: out<=0;
   39634: out<=1;
   39635: out<=1;
   39636: out<=1;
   39637: out<=0;
   39638: out<=1;
   39639: out<=0;
   39640: out<=0;
   39641: out<=1;
   39642: out<=1;
   39643: out<=0;
   39644: out<=1;
   39645: out<=1;
   39646: out<=1;
   39647: out<=1;
   39648: out<=1;
   39649: out<=1;
   39650: out<=1;
   39651: out<=1;
   39652: out<=0;
   39653: out<=1;
   39654: out<=1;
   39655: out<=0;
   39656: out<=0;
   39657: out<=1;
   39658: out<=0;
   39659: out<=1;
   39660: out<=1;
   39661: out<=1;
   39662: out<=0;
   39663: out<=0;
   39664: out<=1;
   39665: out<=0;
   39666: out<=0;
   39667: out<=1;
   39668: out<=1;
   39669: out<=1;
   39670: out<=1;
   39671: out<=1;
   39672: out<=1;
   39673: out<=1;
   39674: out<=0;
   39675: out<=0;
   39676: out<=1;
   39677: out<=0;
   39678: out<=1;
   39679: out<=0;
   39680: out<=1;
   39681: out<=1;
   39682: out<=0;
   39683: out<=0;
   39684: out<=0;
   39685: out<=1;
   39686: out<=0;
   39687: out<=1;
   39688: out<=1;
   39689: out<=0;
   39690: out<=0;
   39691: out<=1;
   39692: out<=0;
   39693: out<=0;
   39694: out<=0;
   39695: out<=0;
   39696: out<=0;
   39697: out<=1;
   39698: out<=0;
   39699: out<=1;
   39700: out<=0;
   39701: out<=0;
   39702: out<=1;
   39703: out<=1;
   39704: out<=1;
   39705: out<=1;
   39706: out<=1;
   39707: out<=1;
   39708: out<=1;
   39709: out<=0;
   39710: out<=0;
   39711: out<=1;
   39712: out<=0;
   39713: out<=1;
   39714: out<=1;
   39715: out<=0;
   39716: out<=0;
   39717: out<=0;
   39718: out<=0;
   39719: out<=0;
   39720: out<=0;
   39721: out<=0;
   39722: out<=1;
   39723: out<=1;
   39724: out<=0;
   39725: out<=1;
   39726: out<=0;
   39727: out<=1;
   39728: out<=1;
   39729: out<=1;
   39730: out<=1;
   39731: out<=1;
   39732: out<=0;
   39733: out<=1;
   39734: out<=1;
   39735: out<=0;
   39736: out<=0;
   39737: out<=1;
   39738: out<=0;
   39739: out<=1;
   39740: out<=1;
   39741: out<=1;
   39742: out<=0;
   39743: out<=0;
   39744: out<=0;
   39745: out<=0;
   39746: out<=1;
   39747: out<=1;
   39748: out<=1;
   39749: out<=0;
   39750: out<=1;
   39751: out<=0;
   39752: out<=0;
   39753: out<=1;
   39754: out<=1;
   39755: out<=0;
   39756: out<=1;
   39757: out<=1;
   39758: out<=1;
   39759: out<=1;
   39760: out<=0;
   39761: out<=1;
   39762: out<=0;
   39763: out<=1;
   39764: out<=0;
   39765: out<=0;
   39766: out<=1;
   39767: out<=1;
   39768: out<=1;
   39769: out<=1;
   39770: out<=1;
   39771: out<=1;
   39772: out<=1;
   39773: out<=0;
   39774: out<=0;
   39775: out<=1;
   39776: out<=0;
   39777: out<=1;
   39778: out<=1;
   39779: out<=0;
   39780: out<=0;
   39781: out<=0;
   39782: out<=0;
   39783: out<=0;
   39784: out<=0;
   39785: out<=0;
   39786: out<=1;
   39787: out<=1;
   39788: out<=0;
   39789: out<=1;
   39790: out<=0;
   39791: out<=1;
   39792: out<=0;
   39793: out<=0;
   39794: out<=0;
   39795: out<=0;
   39796: out<=1;
   39797: out<=0;
   39798: out<=0;
   39799: out<=1;
   39800: out<=1;
   39801: out<=0;
   39802: out<=1;
   39803: out<=0;
   39804: out<=0;
   39805: out<=0;
   39806: out<=1;
   39807: out<=1;
   39808: out<=0;
   39809: out<=0;
   39810: out<=1;
   39811: out<=1;
   39812: out<=1;
   39813: out<=0;
   39814: out<=1;
   39815: out<=0;
   39816: out<=0;
   39817: out<=1;
   39818: out<=1;
   39819: out<=0;
   39820: out<=1;
   39821: out<=1;
   39822: out<=1;
   39823: out<=1;
   39824: out<=0;
   39825: out<=1;
   39826: out<=0;
   39827: out<=1;
   39828: out<=0;
   39829: out<=0;
   39830: out<=1;
   39831: out<=1;
   39832: out<=1;
   39833: out<=1;
   39834: out<=1;
   39835: out<=1;
   39836: out<=1;
   39837: out<=0;
   39838: out<=0;
   39839: out<=1;
   39840: out<=1;
   39841: out<=0;
   39842: out<=0;
   39843: out<=1;
   39844: out<=1;
   39845: out<=1;
   39846: out<=1;
   39847: out<=1;
   39848: out<=1;
   39849: out<=1;
   39850: out<=0;
   39851: out<=0;
   39852: out<=1;
   39853: out<=0;
   39854: out<=1;
   39855: out<=0;
   39856: out<=1;
   39857: out<=1;
   39858: out<=1;
   39859: out<=1;
   39860: out<=0;
   39861: out<=1;
   39862: out<=1;
   39863: out<=0;
   39864: out<=0;
   39865: out<=1;
   39866: out<=0;
   39867: out<=1;
   39868: out<=1;
   39869: out<=1;
   39870: out<=0;
   39871: out<=0;
   39872: out<=1;
   39873: out<=1;
   39874: out<=0;
   39875: out<=0;
   39876: out<=0;
   39877: out<=1;
   39878: out<=0;
   39879: out<=1;
   39880: out<=1;
   39881: out<=0;
   39882: out<=0;
   39883: out<=1;
   39884: out<=0;
   39885: out<=0;
   39886: out<=0;
   39887: out<=0;
   39888: out<=0;
   39889: out<=1;
   39890: out<=0;
   39891: out<=1;
   39892: out<=0;
   39893: out<=0;
   39894: out<=1;
   39895: out<=1;
   39896: out<=1;
   39897: out<=1;
   39898: out<=1;
   39899: out<=1;
   39900: out<=1;
   39901: out<=0;
   39902: out<=0;
   39903: out<=1;
   39904: out<=1;
   39905: out<=0;
   39906: out<=0;
   39907: out<=1;
   39908: out<=1;
   39909: out<=1;
   39910: out<=1;
   39911: out<=1;
   39912: out<=1;
   39913: out<=1;
   39914: out<=0;
   39915: out<=0;
   39916: out<=1;
   39917: out<=0;
   39918: out<=1;
   39919: out<=0;
   39920: out<=0;
   39921: out<=0;
   39922: out<=0;
   39923: out<=0;
   39924: out<=1;
   39925: out<=0;
   39926: out<=0;
   39927: out<=1;
   39928: out<=1;
   39929: out<=0;
   39930: out<=1;
   39931: out<=0;
   39932: out<=0;
   39933: out<=0;
   39934: out<=1;
   39935: out<=1;
   39936: out<=0;
   39937: out<=1;
   39938: out<=1;
   39939: out<=0;
   39940: out<=1;
   39941: out<=1;
   39942: out<=1;
   39943: out<=1;
   39944: out<=1;
   39945: out<=1;
   39946: out<=0;
   39947: out<=0;
   39948: out<=0;
   39949: out<=1;
   39950: out<=0;
   39951: out<=1;
   39952: out<=1;
   39953: out<=1;
   39954: out<=1;
   39955: out<=1;
   39956: out<=1;
   39957: out<=0;
   39958: out<=0;
   39959: out<=1;
   39960: out<=1;
   39961: out<=0;
   39962: out<=1;
   39963: out<=0;
   39964: out<=1;
   39965: out<=1;
   39966: out<=0;
   39967: out<=0;
   39968: out<=0;
   39969: out<=0;
   39970: out<=1;
   39971: out<=1;
   39972: out<=0;
   39973: out<=1;
   39974: out<=0;
   39975: out<=1;
   39976: out<=1;
   39977: out<=0;
   39978: out<=0;
   39979: out<=1;
   39980: out<=1;
   39981: out<=1;
   39982: out<=1;
   39983: out<=1;
   39984: out<=1;
   39985: out<=0;
   39986: out<=1;
   39987: out<=0;
   39988: out<=0;
   39989: out<=0;
   39990: out<=1;
   39991: out<=1;
   39992: out<=1;
   39993: out<=1;
   39994: out<=1;
   39995: out<=1;
   39996: out<=0;
   39997: out<=1;
   39998: out<=1;
   39999: out<=0;
   40000: out<=0;
   40001: out<=1;
   40002: out<=1;
   40003: out<=0;
   40004: out<=1;
   40005: out<=1;
   40006: out<=1;
   40007: out<=1;
   40008: out<=1;
   40009: out<=1;
   40010: out<=0;
   40011: out<=0;
   40012: out<=0;
   40013: out<=1;
   40014: out<=0;
   40015: out<=1;
   40016: out<=0;
   40017: out<=0;
   40018: out<=0;
   40019: out<=0;
   40020: out<=0;
   40021: out<=1;
   40022: out<=1;
   40023: out<=0;
   40024: out<=0;
   40025: out<=1;
   40026: out<=0;
   40027: out<=1;
   40028: out<=0;
   40029: out<=0;
   40030: out<=1;
   40031: out<=1;
   40032: out<=1;
   40033: out<=1;
   40034: out<=0;
   40035: out<=0;
   40036: out<=1;
   40037: out<=0;
   40038: out<=1;
   40039: out<=0;
   40040: out<=0;
   40041: out<=1;
   40042: out<=1;
   40043: out<=0;
   40044: out<=0;
   40045: out<=0;
   40046: out<=0;
   40047: out<=0;
   40048: out<=1;
   40049: out<=0;
   40050: out<=1;
   40051: out<=0;
   40052: out<=0;
   40053: out<=0;
   40054: out<=1;
   40055: out<=1;
   40056: out<=1;
   40057: out<=1;
   40058: out<=1;
   40059: out<=1;
   40060: out<=0;
   40061: out<=1;
   40062: out<=1;
   40063: out<=0;
   40064: out<=1;
   40065: out<=0;
   40066: out<=0;
   40067: out<=1;
   40068: out<=0;
   40069: out<=0;
   40070: out<=0;
   40071: out<=0;
   40072: out<=0;
   40073: out<=0;
   40074: out<=1;
   40075: out<=1;
   40076: out<=1;
   40077: out<=0;
   40078: out<=1;
   40079: out<=0;
   40080: out<=1;
   40081: out<=1;
   40082: out<=1;
   40083: out<=1;
   40084: out<=1;
   40085: out<=0;
   40086: out<=0;
   40087: out<=1;
   40088: out<=1;
   40089: out<=0;
   40090: out<=1;
   40091: out<=0;
   40092: out<=1;
   40093: out<=1;
   40094: out<=0;
   40095: out<=0;
   40096: out<=1;
   40097: out<=1;
   40098: out<=0;
   40099: out<=0;
   40100: out<=1;
   40101: out<=0;
   40102: out<=1;
   40103: out<=0;
   40104: out<=0;
   40105: out<=1;
   40106: out<=1;
   40107: out<=0;
   40108: out<=0;
   40109: out<=0;
   40110: out<=0;
   40111: out<=0;
   40112: out<=1;
   40113: out<=0;
   40114: out<=1;
   40115: out<=0;
   40116: out<=0;
   40117: out<=0;
   40118: out<=1;
   40119: out<=1;
   40120: out<=1;
   40121: out<=1;
   40122: out<=1;
   40123: out<=1;
   40124: out<=0;
   40125: out<=1;
   40126: out<=1;
   40127: out<=0;
   40128: out<=1;
   40129: out<=0;
   40130: out<=0;
   40131: out<=1;
   40132: out<=0;
   40133: out<=0;
   40134: out<=0;
   40135: out<=0;
   40136: out<=0;
   40137: out<=0;
   40138: out<=1;
   40139: out<=1;
   40140: out<=1;
   40141: out<=0;
   40142: out<=1;
   40143: out<=0;
   40144: out<=0;
   40145: out<=0;
   40146: out<=0;
   40147: out<=0;
   40148: out<=0;
   40149: out<=1;
   40150: out<=1;
   40151: out<=0;
   40152: out<=0;
   40153: out<=1;
   40154: out<=0;
   40155: out<=1;
   40156: out<=0;
   40157: out<=0;
   40158: out<=1;
   40159: out<=1;
   40160: out<=0;
   40161: out<=0;
   40162: out<=1;
   40163: out<=1;
   40164: out<=0;
   40165: out<=1;
   40166: out<=0;
   40167: out<=1;
   40168: out<=1;
   40169: out<=0;
   40170: out<=0;
   40171: out<=1;
   40172: out<=1;
   40173: out<=1;
   40174: out<=1;
   40175: out<=1;
   40176: out<=1;
   40177: out<=0;
   40178: out<=1;
   40179: out<=0;
   40180: out<=0;
   40181: out<=0;
   40182: out<=1;
   40183: out<=1;
   40184: out<=1;
   40185: out<=1;
   40186: out<=1;
   40187: out<=1;
   40188: out<=0;
   40189: out<=1;
   40190: out<=1;
   40191: out<=0;
   40192: out<=0;
   40193: out<=0;
   40194: out<=0;
   40195: out<=0;
   40196: out<=0;
   40197: out<=1;
   40198: out<=1;
   40199: out<=0;
   40200: out<=0;
   40201: out<=1;
   40202: out<=0;
   40203: out<=1;
   40204: out<=0;
   40205: out<=0;
   40206: out<=1;
   40207: out<=1;
   40208: out<=0;
   40209: out<=1;
   40210: out<=1;
   40211: out<=0;
   40212: out<=1;
   40213: out<=1;
   40214: out<=1;
   40215: out<=1;
   40216: out<=1;
   40217: out<=1;
   40218: out<=0;
   40219: out<=0;
   40220: out<=0;
   40221: out<=1;
   40222: out<=0;
   40223: out<=1;
   40224: out<=1;
   40225: out<=0;
   40226: out<=1;
   40227: out<=0;
   40228: out<=0;
   40229: out<=0;
   40230: out<=1;
   40231: out<=1;
   40232: out<=1;
   40233: out<=1;
   40234: out<=1;
   40235: out<=1;
   40236: out<=0;
   40237: out<=1;
   40238: out<=1;
   40239: out<=0;
   40240: out<=1;
   40241: out<=1;
   40242: out<=0;
   40243: out<=0;
   40244: out<=1;
   40245: out<=0;
   40246: out<=1;
   40247: out<=0;
   40248: out<=0;
   40249: out<=1;
   40250: out<=1;
   40251: out<=0;
   40252: out<=0;
   40253: out<=0;
   40254: out<=0;
   40255: out<=0;
   40256: out<=1;
   40257: out<=1;
   40258: out<=1;
   40259: out<=1;
   40260: out<=1;
   40261: out<=0;
   40262: out<=0;
   40263: out<=1;
   40264: out<=1;
   40265: out<=0;
   40266: out<=1;
   40267: out<=0;
   40268: out<=1;
   40269: out<=1;
   40270: out<=0;
   40271: out<=0;
   40272: out<=0;
   40273: out<=1;
   40274: out<=1;
   40275: out<=0;
   40276: out<=1;
   40277: out<=1;
   40278: out<=1;
   40279: out<=1;
   40280: out<=1;
   40281: out<=1;
   40282: out<=0;
   40283: out<=0;
   40284: out<=0;
   40285: out<=1;
   40286: out<=0;
   40287: out<=1;
   40288: out<=1;
   40289: out<=0;
   40290: out<=1;
   40291: out<=0;
   40292: out<=0;
   40293: out<=0;
   40294: out<=1;
   40295: out<=1;
   40296: out<=1;
   40297: out<=1;
   40298: out<=1;
   40299: out<=1;
   40300: out<=0;
   40301: out<=1;
   40302: out<=1;
   40303: out<=0;
   40304: out<=0;
   40305: out<=0;
   40306: out<=1;
   40307: out<=1;
   40308: out<=0;
   40309: out<=1;
   40310: out<=0;
   40311: out<=1;
   40312: out<=1;
   40313: out<=0;
   40314: out<=0;
   40315: out<=1;
   40316: out<=1;
   40317: out<=1;
   40318: out<=1;
   40319: out<=1;
   40320: out<=0;
   40321: out<=0;
   40322: out<=0;
   40323: out<=0;
   40324: out<=0;
   40325: out<=1;
   40326: out<=1;
   40327: out<=0;
   40328: out<=0;
   40329: out<=1;
   40330: out<=0;
   40331: out<=1;
   40332: out<=0;
   40333: out<=0;
   40334: out<=1;
   40335: out<=1;
   40336: out<=1;
   40337: out<=0;
   40338: out<=0;
   40339: out<=1;
   40340: out<=0;
   40341: out<=0;
   40342: out<=0;
   40343: out<=0;
   40344: out<=0;
   40345: out<=0;
   40346: out<=1;
   40347: out<=1;
   40348: out<=1;
   40349: out<=0;
   40350: out<=1;
   40351: out<=0;
   40352: out<=1;
   40353: out<=0;
   40354: out<=1;
   40355: out<=0;
   40356: out<=0;
   40357: out<=0;
   40358: out<=1;
   40359: out<=1;
   40360: out<=1;
   40361: out<=1;
   40362: out<=1;
   40363: out<=1;
   40364: out<=0;
   40365: out<=1;
   40366: out<=1;
   40367: out<=0;
   40368: out<=0;
   40369: out<=0;
   40370: out<=1;
   40371: out<=1;
   40372: out<=0;
   40373: out<=1;
   40374: out<=0;
   40375: out<=1;
   40376: out<=1;
   40377: out<=0;
   40378: out<=0;
   40379: out<=1;
   40380: out<=1;
   40381: out<=1;
   40382: out<=1;
   40383: out<=1;
   40384: out<=1;
   40385: out<=1;
   40386: out<=1;
   40387: out<=1;
   40388: out<=1;
   40389: out<=0;
   40390: out<=0;
   40391: out<=1;
   40392: out<=1;
   40393: out<=0;
   40394: out<=1;
   40395: out<=0;
   40396: out<=1;
   40397: out<=1;
   40398: out<=0;
   40399: out<=0;
   40400: out<=1;
   40401: out<=0;
   40402: out<=0;
   40403: out<=1;
   40404: out<=0;
   40405: out<=0;
   40406: out<=0;
   40407: out<=0;
   40408: out<=0;
   40409: out<=0;
   40410: out<=1;
   40411: out<=1;
   40412: out<=1;
   40413: out<=0;
   40414: out<=1;
   40415: out<=0;
   40416: out<=1;
   40417: out<=0;
   40418: out<=1;
   40419: out<=0;
   40420: out<=0;
   40421: out<=0;
   40422: out<=1;
   40423: out<=1;
   40424: out<=1;
   40425: out<=1;
   40426: out<=1;
   40427: out<=1;
   40428: out<=0;
   40429: out<=1;
   40430: out<=1;
   40431: out<=0;
   40432: out<=1;
   40433: out<=1;
   40434: out<=0;
   40435: out<=0;
   40436: out<=1;
   40437: out<=0;
   40438: out<=1;
   40439: out<=0;
   40440: out<=0;
   40441: out<=1;
   40442: out<=1;
   40443: out<=0;
   40444: out<=0;
   40445: out<=0;
   40446: out<=0;
   40447: out<=0;
   40448: out<=1;
   40449: out<=1;
   40450: out<=0;
   40451: out<=0;
   40452: out<=1;
   40453: out<=0;
   40454: out<=1;
   40455: out<=0;
   40456: out<=0;
   40457: out<=1;
   40458: out<=1;
   40459: out<=0;
   40460: out<=0;
   40461: out<=0;
   40462: out<=0;
   40463: out<=0;
   40464: out<=1;
   40465: out<=0;
   40466: out<=1;
   40467: out<=0;
   40468: out<=0;
   40469: out<=0;
   40470: out<=1;
   40471: out<=1;
   40472: out<=1;
   40473: out<=1;
   40474: out<=1;
   40475: out<=1;
   40476: out<=0;
   40477: out<=1;
   40478: out<=1;
   40479: out<=0;
   40480: out<=1;
   40481: out<=0;
   40482: out<=0;
   40483: out<=1;
   40484: out<=0;
   40485: out<=0;
   40486: out<=0;
   40487: out<=0;
   40488: out<=0;
   40489: out<=0;
   40490: out<=1;
   40491: out<=1;
   40492: out<=1;
   40493: out<=0;
   40494: out<=1;
   40495: out<=0;
   40496: out<=1;
   40497: out<=1;
   40498: out<=1;
   40499: out<=1;
   40500: out<=1;
   40501: out<=0;
   40502: out<=0;
   40503: out<=1;
   40504: out<=1;
   40505: out<=0;
   40506: out<=1;
   40507: out<=0;
   40508: out<=1;
   40509: out<=1;
   40510: out<=0;
   40511: out<=0;
   40512: out<=0;
   40513: out<=0;
   40514: out<=1;
   40515: out<=1;
   40516: out<=0;
   40517: out<=1;
   40518: out<=0;
   40519: out<=1;
   40520: out<=1;
   40521: out<=0;
   40522: out<=0;
   40523: out<=1;
   40524: out<=1;
   40525: out<=1;
   40526: out<=1;
   40527: out<=1;
   40528: out<=1;
   40529: out<=0;
   40530: out<=1;
   40531: out<=0;
   40532: out<=0;
   40533: out<=0;
   40534: out<=1;
   40535: out<=1;
   40536: out<=1;
   40537: out<=1;
   40538: out<=1;
   40539: out<=1;
   40540: out<=0;
   40541: out<=1;
   40542: out<=1;
   40543: out<=0;
   40544: out<=1;
   40545: out<=0;
   40546: out<=0;
   40547: out<=1;
   40548: out<=0;
   40549: out<=0;
   40550: out<=0;
   40551: out<=0;
   40552: out<=0;
   40553: out<=0;
   40554: out<=1;
   40555: out<=1;
   40556: out<=1;
   40557: out<=0;
   40558: out<=1;
   40559: out<=0;
   40560: out<=0;
   40561: out<=0;
   40562: out<=0;
   40563: out<=0;
   40564: out<=0;
   40565: out<=1;
   40566: out<=1;
   40567: out<=0;
   40568: out<=0;
   40569: out<=1;
   40570: out<=0;
   40571: out<=1;
   40572: out<=0;
   40573: out<=0;
   40574: out<=1;
   40575: out<=1;
   40576: out<=0;
   40577: out<=0;
   40578: out<=1;
   40579: out<=1;
   40580: out<=0;
   40581: out<=1;
   40582: out<=0;
   40583: out<=1;
   40584: out<=1;
   40585: out<=0;
   40586: out<=0;
   40587: out<=1;
   40588: out<=1;
   40589: out<=1;
   40590: out<=1;
   40591: out<=1;
   40592: out<=1;
   40593: out<=0;
   40594: out<=1;
   40595: out<=0;
   40596: out<=0;
   40597: out<=0;
   40598: out<=1;
   40599: out<=1;
   40600: out<=1;
   40601: out<=1;
   40602: out<=1;
   40603: out<=1;
   40604: out<=0;
   40605: out<=1;
   40606: out<=1;
   40607: out<=0;
   40608: out<=0;
   40609: out<=1;
   40610: out<=1;
   40611: out<=0;
   40612: out<=1;
   40613: out<=1;
   40614: out<=1;
   40615: out<=1;
   40616: out<=1;
   40617: out<=1;
   40618: out<=0;
   40619: out<=0;
   40620: out<=0;
   40621: out<=1;
   40622: out<=0;
   40623: out<=1;
   40624: out<=1;
   40625: out<=1;
   40626: out<=1;
   40627: out<=1;
   40628: out<=1;
   40629: out<=0;
   40630: out<=0;
   40631: out<=1;
   40632: out<=1;
   40633: out<=0;
   40634: out<=1;
   40635: out<=0;
   40636: out<=1;
   40637: out<=1;
   40638: out<=0;
   40639: out<=0;
   40640: out<=1;
   40641: out<=1;
   40642: out<=0;
   40643: out<=0;
   40644: out<=1;
   40645: out<=0;
   40646: out<=1;
   40647: out<=0;
   40648: out<=0;
   40649: out<=1;
   40650: out<=1;
   40651: out<=0;
   40652: out<=0;
   40653: out<=0;
   40654: out<=0;
   40655: out<=0;
   40656: out<=1;
   40657: out<=0;
   40658: out<=1;
   40659: out<=0;
   40660: out<=0;
   40661: out<=0;
   40662: out<=1;
   40663: out<=1;
   40664: out<=1;
   40665: out<=1;
   40666: out<=1;
   40667: out<=1;
   40668: out<=0;
   40669: out<=1;
   40670: out<=1;
   40671: out<=0;
   40672: out<=0;
   40673: out<=1;
   40674: out<=1;
   40675: out<=0;
   40676: out<=1;
   40677: out<=1;
   40678: out<=1;
   40679: out<=1;
   40680: out<=1;
   40681: out<=1;
   40682: out<=0;
   40683: out<=0;
   40684: out<=0;
   40685: out<=1;
   40686: out<=0;
   40687: out<=1;
   40688: out<=0;
   40689: out<=0;
   40690: out<=0;
   40691: out<=0;
   40692: out<=0;
   40693: out<=1;
   40694: out<=1;
   40695: out<=0;
   40696: out<=0;
   40697: out<=1;
   40698: out<=0;
   40699: out<=1;
   40700: out<=0;
   40701: out<=0;
   40702: out<=1;
   40703: out<=1;
   40704: out<=1;
   40705: out<=0;
   40706: out<=1;
   40707: out<=0;
   40708: out<=0;
   40709: out<=0;
   40710: out<=1;
   40711: out<=1;
   40712: out<=1;
   40713: out<=1;
   40714: out<=1;
   40715: out<=1;
   40716: out<=0;
   40717: out<=1;
   40718: out<=1;
   40719: out<=0;
   40720: out<=0;
   40721: out<=0;
   40722: out<=1;
   40723: out<=1;
   40724: out<=0;
   40725: out<=1;
   40726: out<=0;
   40727: out<=1;
   40728: out<=1;
   40729: out<=0;
   40730: out<=0;
   40731: out<=1;
   40732: out<=1;
   40733: out<=1;
   40734: out<=1;
   40735: out<=1;
   40736: out<=0;
   40737: out<=0;
   40738: out<=0;
   40739: out<=0;
   40740: out<=0;
   40741: out<=1;
   40742: out<=1;
   40743: out<=0;
   40744: out<=0;
   40745: out<=1;
   40746: out<=0;
   40747: out<=1;
   40748: out<=0;
   40749: out<=0;
   40750: out<=1;
   40751: out<=1;
   40752: out<=1;
   40753: out<=0;
   40754: out<=0;
   40755: out<=1;
   40756: out<=0;
   40757: out<=0;
   40758: out<=0;
   40759: out<=0;
   40760: out<=0;
   40761: out<=0;
   40762: out<=1;
   40763: out<=1;
   40764: out<=1;
   40765: out<=0;
   40766: out<=1;
   40767: out<=0;
   40768: out<=1;
   40769: out<=0;
   40770: out<=1;
   40771: out<=0;
   40772: out<=0;
   40773: out<=0;
   40774: out<=1;
   40775: out<=1;
   40776: out<=1;
   40777: out<=1;
   40778: out<=1;
   40779: out<=1;
   40780: out<=0;
   40781: out<=1;
   40782: out<=1;
   40783: out<=0;
   40784: out<=1;
   40785: out<=1;
   40786: out<=0;
   40787: out<=0;
   40788: out<=1;
   40789: out<=0;
   40790: out<=1;
   40791: out<=0;
   40792: out<=0;
   40793: out<=1;
   40794: out<=1;
   40795: out<=0;
   40796: out<=0;
   40797: out<=0;
   40798: out<=0;
   40799: out<=0;
   40800: out<=1;
   40801: out<=1;
   40802: out<=1;
   40803: out<=1;
   40804: out<=1;
   40805: out<=0;
   40806: out<=0;
   40807: out<=1;
   40808: out<=1;
   40809: out<=0;
   40810: out<=1;
   40811: out<=0;
   40812: out<=1;
   40813: out<=1;
   40814: out<=0;
   40815: out<=0;
   40816: out<=1;
   40817: out<=0;
   40818: out<=0;
   40819: out<=1;
   40820: out<=0;
   40821: out<=0;
   40822: out<=0;
   40823: out<=0;
   40824: out<=0;
   40825: out<=0;
   40826: out<=1;
   40827: out<=1;
   40828: out<=1;
   40829: out<=0;
   40830: out<=1;
   40831: out<=0;
   40832: out<=1;
   40833: out<=0;
   40834: out<=1;
   40835: out<=0;
   40836: out<=0;
   40837: out<=0;
   40838: out<=1;
   40839: out<=1;
   40840: out<=1;
   40841: out<=1;
   40842: out<=1;
   40843: out<=1;
   40844: out<=0;
   40845: out<=1;
   40846: out<=1;
   40847: out<=0;
   40848: out<=1;
   40849: out<=1;
   40850: out<=0;
   40851: out<=0;
   40852: out<=1;
   40853: out<=0;
   40854: out<=1;
   40855: out<=0;
   40856: out<=0;
   40857: out<=1;
   40858: out<=1;
   40859: out<=0;
   40860: out<=0;
   40861: out<=0;
   40862: out<=0;
   40863: out<=0;
   40864: out<=0;
   40865: out<=0;
   40866: out<=0;
   40867: out<=0;
   40868: out<=0;
   40869: out<=1;
   40870: out<=1;
   40871: out<=0;
   40872: out<=0;
   40873: out<=1;
   40874: out<=0;
   40875: out<=1;
   40876: out<=0;
   40877: out<=0;
   40878: out<=1;
   40879: out<=1;
   40880: out<=0;
   40881: out<=1;
   40882: out<=1;
   40883: out<=0;
   40884: out<=1;
   40885: out<=1;
   40886: out<=1;
   40887: out<=1;
   40888: out<=1;
   40889: out<=1;
   40890: out<=0;
   40891: out<=0;
   40892: out<=0;
   40893: out<=1;
   40894: out<=0;
   40895: out<=1;
   40896: out<=1;
   40897: out<=0;
   40898: out<=1;
   40899: out<=0;
   40900: out<=0;
   40901: out<=0;
   40902: out<=1;
   40903: out<=1;
   40904: out<=1;
   40905: out<=1;
   40906: out<=1;
   40907: out<=1;
   40908: out<=0;
   40909: out<=1;
   40910: out<=1;
   40911: out<=0;
   40912: out<=0;
   40913: out<=0;
   40914: out<=1;
   40915: out<=1;
   40916: out<=0;
   40917: out<=1;
   40918: out<=0;
   40919: out<=1;
   40920: out<=1;
   40921: out<=0;
   40922: out<=0;
   40923: out<=1;
   40924: out<=1;
   40925: out<=1;
   40926: out<=1;
   40927: out<=1;
   40928: out<=1;
   40929: out<=1;
   40930: out<=1;
   40931: out<=1;
   40932: out<=1;
   40933: out<=0;
   40934: out<=0;
   40935: out<=1;
   40936: out<=1;
   40937: out<=0;
   40938: out<=1;
   40939: out<=0;
   40940: out<=1;
   40941: out<=1;
   40942: out<=0;
   40943: out<=0;
   40944: out<=0;
   40945: out<=1;
   40946: out<=1;
   40947: out<=0;
   40948: out<=1;
   40949: out<=1;
   40950: out<=1;
   40951: out<=1;
   40952: out<=1;
   40953: out<=1;
   40954: out<=0;
   40955: out<=0;
   40956: out<=0;
   40957: out<=1;
   40958: out<=0;
   40959: out<=1;
   40960: out<=0;
   40961: out<=1;
   40962: out<=0;
   40963: out<=1;
   40964: out<=1;
   40965: out<=1;
   40966: out<=0;
   40967: out<=0;
   40968: out<=0;
   40969: out<=0;
   40970: out<=0;
   40971: out<=0;
   40972: out<=1;
   40973: out<=0;
   40974: out<=0;
   40975: out<=1;
   40976: out<=1;
   40977: out<=1;
   40978: out<=0;
   40979: out<=0;
   40980: out<=1;
   40981: out<=0;
   40982: out<=1;
   40983: out<=0;
   40984: out<=0;
   40985: out<=1;
   40986: out<=1;
   40987: out<=0;
   40988: out<=0;
   40989: out<=0;
   40990: out<=0;
   40991: out<=0;
   40992: out<=0;
   40993: out<=0;
   40994: out<=0;
   40995: out<=0;
   40996: out<=0;
   40997: out<=1;
   40998: out<=1;
   40999: out<=0;
   41000: out<=0;
   41001: out<=1;
   41002: out<=0;
   41003: out<=1;
   41004: out<=0;
   41005: out<=0;
   41006: out<=1;
   41007: out<=1;
   41008: out<=1;
   41009: out<=0;
   41010: out<=0;
   41011: out<=1;
   41012: out<=0;
   41013: out<=0;
   41014: out<=0;
   41015: out<=0;
   41016: out<=0;
   41017: out<=0;
   41018: out<=1;
   41019: out<=1;
   41020: out<=1;
   41021: out<=0;
   41022: out<=1;
   41023: out<=0;
   41024: out<=0;
   41025: out<=1;
   41026: out<=0;
   41027: out<=1;
   41028: out<=1;
   41029: out<=1;
   41030: out<=0;
   41031: out<=0;
   41032: out<=0;
   41033: out<=0;
   41034: out<=0;
   41035: out<=0;
   41036: out<=1;
   41037: out<=0;
   41038: out<=0;
   41039: out<=1;
   41040: out<=0;
   41041: out<=0;
   41042: out<=1;
   41043: out<=1;
   41044: out<=0;
   41045: out<=1;
   41046: out<=0;
   41047: out<=1;
   41048: out<=1;
   41049: out<=0;
   41050: out<=0;
   41051: out<=1;
   41052: out<=1;
   41053: out<=1;
   41054: out<=1;
   41055: out<=1;
   41056: out<=1;
   41057: out<=1;
   41058: out<=1;
   41059: out<=1;
   41060: out<=1;
   41061: out<=0;
   41062: out<=0;
   41063: out<=1;
   41064: out<=1;
   41065: out<=0;
   41066: out<=1;
   41067: out<=0;
   41068: out<=1;
   41069: out<=1;
   41070: out<=0;
   41071: out<=0;
   41072: out<=1;
   41073: out<=0;
   41074: out<=0;
   41075: out<=1;
   41076: out<=0;
   41077: out<=0;
   41078: out<=0;
   41079: out<=0;
   41080: out<=0;
   41081: out<=0;
   41082: out<=1;
   41083: out<=1;
   41084: out<=1;
   41085: out<=0;
   41086: out<=1;
   41087: out<=0;
   41088: out<=0;
   41089: out<=1;
   41090: out<=0;
   41091: out<=1;
   41092: out<=1;
   41093: out<=1;
   41094: out<=0;
   41095: out<=0;
   41096: out<=0;
   41097: out<=0;
   41098: out<=0;
   41099: out<=0;
   41100: out<=1;
   41101: out<=0;
   41102: out<=0;
   41103: out<=1;
   41104: out<=0;
   41105: out<=0;
   41106: out<=1;
   41107: out<=1;
   41108: out<=0;
   41109: out<=1;
   41110: out<=0;
   41111: out<=1;
   41112: out<=1;
   41113: out<=0;
   41114: out<=0;
   41115: out<=1;
   41116: out<=1;
   41117: out<=1;
   41118: out<=1;
   41119: out<=1;
   41120: out<=0;
   41121: out<=0;
   41122: out<=0;
   41123: out<=0;
   41124: out<=0;
   41125: out<=1;
   41126: out<=1;
   41127: out<=0;
   41128: out<=0;
   41129: out<=1;
   41130: out<=0;
   41131: out<=1;
   41132: out<=0;
   41133: out<=0;
   41134: out<=1;
   41135: out<=1;
   41136: out<=0;
   41137: out<=1;
   41138: out<=1;
   41139: out<=0;
   41140: out<=1;
   41141: out<=1;
   41142: out<=1;
   41143: out<=1;
   41144: out<=1;
   41145: out<=1;
   41146: out<=0;
   41147: out<=0;
   41148: out<=0;
   41149: out<=1;
   41150: out<=0;
   41151: out<=1;
   41152: out<=0;
   41153: out<=1;
   41154: out<=0;
   41155: out<=1;
   41156: out<=1;
   41157: out<=1;
   41158: out<=0;
   41159: out<=0;
   41160: out<=0;
   41161: out<=0;
   41162: out<=0;
   41163: out<=0;
   41164: out<=1;
   41165: out<=0;
   41166: out<=0;
   41167: out<=1;
   41168: out<=1;
   41169: out<=1;
   41170: out<=0;
   41171: out<=0;
   41172: out<=1;
   41173: out<=0;
   41174: out<=1;
   41175: out<=0;
   41176: out<=0;
   41177: out<=1;
   41178: out<=1;
   41179: out<=0;
   41180: out<=0;
   41181: out<=0;
   41182: out<=0;
   41183: out<=0;
   41184: out<=1;
   41185: out<=1;
   41186: out<=1;
   41187: out<=1;
   41188: out<=1;
   41189: out<=0;
   41190: out<=0;
   41191: out<=1;
   41192: out<=1;
   41193: out<=0;
   41194: out<=1;
   41195: out<=0;
   41196: out<=1;
   41197: out<=1;
   41198: out<=0;
   41199: out<=0;
   41200: out<=0;
   41201: out<=1;
   41202: out<=1;
   41203: out<=0;
   41204: out<=1;
   41205: out<=1;
   41206: out<=1;
   41207: out<=1;
   41208: out<=1;
   41209: out<=1;
   41210: out<=0;
   41211: out<=0;
   41212: out<=0;
   41213: out<=1;
   41214: out<=0;
   41215: out<=1;
   41216: out<=0;
   41217: out<=0;
   41218: out<=1;
   41219: out<=1;
   41220: out<=0;
   41221: out<=1;
   41222: out<=0;
   41223: out<=1;
   41224: out<=1;
   41225: out<=0;
   41226: out<=0;
   41227: out<=1;
   41228: out<=1;
   41229: out<=1;
   41230: out<=1;
   41231: out<=1;
   41232: out<=0;
   41233: out<=1;
   41234: out<=0;
   41235: out<=1;
   41236: out<=1;
   41237: out<=1;
   41238: out<=0;
   41239: out<=0;
   41240: out<=0;
   41241: out<=0;
   41242: out<=0;
   41243: out<=0;
   41244: out<=1;
   41245: out<=0;
   41246: out<=0;
   41247: out<=1;
   41248: out<=1;
   41249: out<=0;
   41250: out<=0;
   41251: out<=1;
   41252: out<=0;
   41253: out<=0;
   41254: out<=0;
   41255: out<=0;
   41256: out<=0;
   41257: out<=0;
   41258: out<=1;
   41259: out<=1;
   41260: out<=1;
   41261: out<=0;
   41262: out<=1;
   41263: out<=0;
   41264: out<=1;
   41265: out<=1;
   41266: out<=1;
   41267: out<=1;
   41268: out<=1;
   41269: out<=0;
   41270: out<=0;
   41271: out<=1;
   41272: out<=1;
   41273: out<=0;
   41274: out<=1;
   41275: out<=0;
   41276: out<=1;
   41277: out<=1;
   41278: out<=0;
   41279: out<=0;
   41280: out<=1;
   41281: out<=1;
   41282: out<=0;
   41283: out<=0;
   41284: out<=1;
   41285: out<=0;
   41286: out<=1;
   41287: out<=0;
   41288: out<=0;
   41289: out<=1;
   41290: out<=1;
   41291: out<=0;
   41292: out<=0;
   41293: out<=0;
   41294: out<=0;
   41295: out<=0;
   41296: out<=0;
   41297: out<=1;
   41298: out<=0;
   41299: out<=1;
   41300: out<=1;
   41301: out<=1;
   41302: out<=0;
   41303: out<=0;
   41304: out<=0;
   41305: out<=0;
   41306: out<=0;
   41307: out<=0;
   41308: out<=1;
   41309: out<=0;
   41310: out<=0;
   41311: out<=1;
   41312: out<=1;
   41313: out<=0;
   41314: out<=0;
   41315: out<=1;
   41316: out<=0;
   41317: out<=0;
   41318: out<=0;
   41319: out<=0;
   41320: out<=0;
   41321: out<=0;
   41322: out<=1;
   41323: out<=1;
   41324: out<=1;
   41325: out<=0;
   41326: out<=1;
   41327: out<=0;
   41328: out<=0;
   41329: out<=0;
   41330: out<=0;
   41331: out<=0;
   41332: out<=0;
   41333: out<=1;
   41334: out<=1;
   41335: out<=0;
   41336: out<=0;
   41337: out<=1;
   41338: out<=0;
   41339: out<=1;
   41340: out<=0;
   41341: out<=0;
   41342: out<=1;
   41343: out<=1;
   41344: out<=1;
   41345: out<=1;
   41346: out<=0;
   41347: out<=0;
   41348: out<=1;
   41349: out<=0;
   41350: out<=1;
   41351: out<=0;
   41352: out<=0;
   41353: out<=1;
   41354: out<=1;
   41355: out<=0;
   41356: out<=0;
   41357: out<=0;
   41358: out<=0;
   41359: out<=0;
   41360: out<=0;
   41361: out<=1;
   41362: out<=0;
   41363: out<=1;
   41364: out<=1;
   41365: out<=1;
   41366: out<=0;
   41367: out<=0;
   41368: out<=0;
   41369: out<=0;
   41370: out<=0;
   41371: out<=0;
   41372: out<=1;
   41373: out<=0;
   41374: out<=0;
   41375: out<=1;
   41376: out<=0;
   41377: out<=1;
   41378: out<=1;
   41379: out<=0;
   41380: out<=1;
   41381: out<=1;
   41382: out<=1;
   41383: out<=1;
   41384: out<=1;
   41385: out<=1;
   41386: out<=0;
   41387: out<=0;
   41388: out<=0;
   41389: out<=1;
   41390: out<=0;
   41391: out<=1;
   41392: out<=1;
   41393: out<=1;
   41394: out<=1;
   41395: out<=1;
   41396: out<=1;
   41397: out<=0;
   41398: out<=0;
   41399: out<=1;
   41400: out<=1;
   41401: out<=0;
   41402: out<=1;
   41403: out<=0;
   41404: out<=1;
   41405: out<=1;
   41406: out<=0;
   41407: out<=0;
   41408: out<=0;
   41409: out<=0;
   41410: out<=1;
   41411: out<=1;
   41412: out<=0;
   41413: out<=1;
   41414: out<=0;
   41415: out<=1;
   41416: out<=1;
   41417: out<=0;
   41418: out<=0;
   41419: out<=1;
   41420: out<=1;
   41421: out<=1;
   41422: out<=1;
   41423: out<=1;
   41424: out<=0;
   41425: out<=1;
   41426: out<=0;
   41427: out<=1;
   41428: out<=1;
   41429: out<=1;
   41430: out<=0;
   41431: out<=0;
   41432: out<=0;
   41433: out<=0;
   41434: out<=0;
   41435: out<=0;
   41436: out<=1;
   41437: out<=0;
   41438: out<=0;
   41439: out<=1;
   41440: out<=0;
   41441: out<=1;
   41442: out<=1;
   41443: out<=0;
   41444: out<=1;
   41445: out<=1;
   41446: out<=1;
   41447: out<=1;
   41448: out<=1;
   41449: out<=1;
   41450: out<=0;
   41451: out<=0;
   41452: out<=0;
   41453: out<=1;
   41454: out<=0;
   41455: out<=1;
   41456: out<=0;
   41457: out<=0;
   41458: out<=0;
   41459: out<=0;
   41460: out<=0;
   41461: out<=1;
   41462: out<=1;
   41463: out<=0;
   41464: out<=0;
   41465: out<=1;
   41466: out<=0;
   41467: out<=1;
   41468: out<=0;
   41469: out<=0;
   41470: out<=1;
   41471: out<=1;
   41472: out<=0;
   41473: out<=0;
   41474: out<=0;
   41475: out<=0;
   41476: out<=0;
   41477: out<=1;
   41478: out<=1;
   41479: out<=0;
   41480: out<=0;
   41481: out<=1;
   41482: out<=0;
   41483: out<=1;
   41484: out<=0;
   41485: out<=0;
   41486: out<=1;
   41487: out<=1;
   41488: out<=0;
   41489: out<=1;
   41490: out<=1;
   41491: out<=0;
   41492: out<=1;
   41493: out<=1;
   41494: out<=1;
   41495: out<=1;
   41496: out<=1;
   41497: out<=1;
   41498: out<=0;
   41499: out<=0;
   41500: out<=0;
   41501: out<=1;
   41502: out<=0;
   41503: out<=1;
   41504: out<=0;
   41505: out<=1;
   41506: out<=0;
   41507: out<=1;
   41508: out<=1;
   41509: out<=1;
   41510: out<=0;
   41511: out<=0;
   41512: out<=0;
   41513: out<=0;
   41514: out<=0;
   41515: out<=0;
   41516: out<=1;
   41517: out<=0;
   41518: out<=0;
   41519: out<=1;
   41520: out<=0;
   41521: out<=0;
   41522: out<=1;
   41523: out<=1;
   41524: out<=0;
   41525: out<=1;
   41526: out<=0;
   41527: out<=1;
   41528: out<=1;
   41529: out<=0;
   41530: out<=0;
   41531: out<=1;
   41532: out<=1;
   41533: out<=1;
   41534: out<=1;
   41535: out<=1;
   41536: out<=1;
   41537: out<=1;
   41538: out<=1;
   41539: out<=1;
   41540: out<=1;
   41541: out<=0;
   41542: out<=0;
   41543: out<=1;
   41544: out<=1;
   41545: out<=0;
   41546: out<=1;
   41547: out<=0;
   41548: out<=1;
   41549: out<=1;
   41550: out<=0;
   41551: out<=0;
   41552: out<=0;
   41553: out<=1;
   41554: out<=1;
   41555: out<=0;
   41556: out<=1;
   41557: out<=1;
   41558: out<=1;
   41559: out<=1;
   41560: out<=1;
   41561: out<=1;
   41562: out<=0;
   41563: out<=0;
   41564: out<=0;
   41565: out<=1;
   41566: out<=0;
   41567: out<=1;
   41568: out<=0;
   41569: out<=1;
   41570: out<=0;
   41571: out<=1;
   41572: out<=1;
   41573: out<=1;
   41574: out<=0;
   41575: out<=0;
   41576: out<=0;
   41577: out<=0;
   41578: out<=0;
   41579: out<=0;
   41580: out<=1;
   41581: out<=0;
   41582: out<=0;
   41583: out<=1;
   41584: out<=1;
   41585: out<=1;
   41586: out<=0;
   41587: out<=0;
   41588: out<=1;
   41589: out<=0;
   41590: out<=1;
   41591: out<=0;
   41592: out<=0;
   41593: out<=1;
   41594: out<=1;
   41595: out<=0;
   41596: out<=0;
   41597: out<=0;
   41598: out<=0;
   41599: out<=0;
   41600: out<=0;
   41601: out<=0;
   41602: out<=0;
   41603: out<=0;
   41604: out<=0;
   41605: out<=1;
   41606: out<=1;
   41607: out<=0;
   41608: out<=0;
   41609: out<=1;
   41610: out<=0;
   41611: out<=1;
   41612: out<=0;
   41613: out<=0;
   41614: out<=1;
   41615: out<=1;
   41616: out<=1;
   41617: out<=0;
   41618: out<=0;
   41619: out<=1;
   41620: out<=0;
   41621: out<=0;
   41622: out<=0;
   41623: out<=0;
   41624: out<=0;
   41625: out<=0;
   41626: out<=1;
   41627: out<=1;
   41628: out<=1;
   41629: out<=0;
   41630: out<=1;
   41631: out<=0;
   41632: out<=0;
   41633: out<=1;
   41634: out<=0;
   41635: out<=1;
   41636: out<=1;
   41637: out<=1;
   41638: out<=0;
   41639: out<=0;
   41640: out<=0;
   41641: out<=0;
   41642: out<=0;
   41643: out<=0;
   41644: out<=1;
   41645: out<=0;
   41646: out<=0;
   41647: out<=1;
   41648: out<=1;
   41649: out<=1;
   41650: out<=0;
   41651: out<=0;
   41652: out<=1;
   41653: out<=0;
   41654: out<=1;
   41655: out<=0;
   41656: out<=0;
   41657: out<=1;
   41658: out<=1;
   41659: out<=0;
   41660: out<=0;
   41661: out<=0;
   41662: out<=0;
   41663: out<=0;
   41664: out<=1;
   41665: out<=1;
   41666: out<=1;
   41667: out<=1;
   41668: out<=1;
   41669: out<=0;
   41670: out<=0;
   41671: out<=1;
   41672: out<=1;
   41673: out<=0;
   41674: out<=1;
   41675: out<=0;
   41676: out<=1;
   41677: out<=1;
   41678: out<=0;
   41679: out<=0;
   41680: out<=1;
   41681: out<=0;
   41682: out<=0;
   41683: out<=1;
   41684: out<=0;
   41685: out<=0;
   41686: out<=0;
   41687: out<=0;
   41688: out<=0;
   41689: out<=0;
   41690: out<=1;
   41691: out<=1;
   41692: out<=1;
   41693: out<=0;
   41694: out<=1;
   41695: out<=0;
   41696: out<=0;
   41697: out<=1;
   41698: out<=0;
   41699: out<=1;
   41700: out<=1;
   41701: out<=1;
   41702: out<=0;
   41703: out<=0;
   41704: out<=0;
   41705: out<=0;
   41706: out<=0;
   41707: out<=0;
   41708: out<=1;
   41709: out<=0;
   41710: out<=0;
   41711: out<=1;
   41712: out<=0;
   41713: out<=0;
   41714: out<=1;
   41715: out<=1;
   41716: out<=0;
   41717: out<=1;
   41718: out<=0;
   41719: out<=1;
   41720: out<=1;
   41721: out<=0;
   41722: out<=0;
   41723: out<=1;
   41724: out<=1;
   41725: out<=1;
   41726: out<=1;
   41727: out<=1;
   41728: out<=0;
   41729: out<=1;
   41730: out<=1;
   41731: out<=0;
   41732: out<=1;
   41733: out<=1;
   41734: out<=1;
   41735: out<=1;
   41736: out<=1;
   41737: out<=1;
   41738: out<=0;
   41739: out<=0;
   41740: out<=0;
   41741: out<=1;
   41742: out<=0;
   41743: out<=1;
   41744: out<=1;
   41745: out<=1;
   41746: out<=1;
   41747: out<=1;
   41748: out<=1;
   41749: out<=0;
   41750: out<=0;
   41751: out<=1;
   41752: out<=1;
   41753: out<=0;
   41754: out<=1;
   41755: out<=0;
   41756: out<=1;
   41757: out<=1;
   41758: out<=0;
   41759: out<=0;
   41760: out<=1;
   41761: out<=1;
   41762: out<=0;
   41763: out<=0;
   41764: out<=1;
   41765: out<=0;
   41766: out<=1;
   41767: out<=0;
   41768: out<=0;
   41769: out<=1;
   41770: out<=1;
   41771: out<=0;
   41772: out<=0;
   41773: out<=0;
   41774: out<=0;
   41775: out<=0;
   41776: out<=0;
   41777: out<=1;
   41778: out<=0;
   41779: out<=1;
   41780: out<=1;
   41781: out<=1;
   41782: out<=0;
   41783: out<=0;
   41784: out<=0;
   41785: out<=0;
   41786: out<=0;
   41787: out<=0;
   41788: out<=1;
   41789: out<=0;
   41790: out<=0;
   41791: out<=1;
   41792: out<=0;
   41793: out<=1;
   41794: out<=1;
   41795: out<=0;
   41796: out<=1;
   41797: out<=1;
   41798: out<=1;
   41799: out<=1;
   41800: out<=1;
   41801: out<=1;
   41802: out<=0;
   41803: out<=0;
   41804: out<=0;
   41805: out<=1;
   41806: out<=0;
   41807: out<=1;
   41808: out<=0;
   41809: out<=0;
   41810: out<=0;
   41811: out<=0;
   41812: out<=0;
   41813: out<=1;
   41814: out<=1;
   41815: out<=0;
   41816: out<=0;
   41817: out<=1;
   41818: out<=0;
   41819: out<=1;
   41820: out<=0;
   41821: out<=0;
   41822: out<=1;
   41823: out<=1;
   41824: out<=0;
   41825: out<=0;
   41826: out<=1;
   41827: out<=1;
   41828: out<=0;
   41829: out<=1;
   41830: out<=0;
   41831: out<=1;
   41832: out<=1;
   41833: out<=0;
   41834: out<=0;
   41835: out<=1;
   41836: out<=1;
   41837: out<=1;
   41838: out<=1;
   41839: out<=1;
   41840: out<=0;
   41841: out<=1;
   41842: out<=0;
   41843: out<=1;
   41844: out<=1;
   41845: out<=1;
   41846: out<=0;
   41847: out<=0;
   41848: out<=0;
   41849: out<=0;
   41850: out<=0;
   41851: out<=0;
   41852: out<=1;
   41853: out<=0;
   41854: out<=0;
   41855: out<=1;
   41856: out<=1;
   41857: out<=0;
   41858: out<=0;
   41859: out<=1;
   41860: out<=0;
   41861: out<=0;
   41862: out<=0;
   41863: out<=0;
   41864: out<=0;
   41865: out<=0;
   41866: out<=1;
   41867: out<=1;
   41868: out<=1;
   41869: out<=0;
   41870: out<=1;
   41871: out<=0;
   41872: out<=1;
   41873: out<=1;
   41874: out<=1;
   41875: out<=1;
   41876: out<=1;
   41877: out<=0;
   41878: out<=0;
   41879: out<=1;
   41880: out<=1;
   41881: out<=0;
   41882: out<=1;
   41883: out<=0;
   41884: out<=1;
   41885: out<=1;
   41886: out<=0;
   41887: out<=0;
   41888: out<=0;
   41889: out<=0;
   41890: out<=1;
   41891: out<=1;
   41892: out<=0;
   41893: out<=1;
   41894: out<=0;
   41895: out<=1;
   41896: out<=1;
   41897: out<=0;
   41898: out<=0;
   41899: out<=1;
   41900: out<=1;
   41901: out<=1;
   41902: out<=1;
   41903: out<=1;
   41904: out<=0;
   41905: out<=1;
   41906: out<=0;
   41907: out<=1;
   41908: out<=1;
   41909: out<=1;
   41910: out<=0;
   41911: out<=0;
   41912: out<=0;
   41913: out<=0;
   41914: out<=0;
   41915: out<=0;
   41916: out<=1;
   41917: out<=0;
   41918: out<=0;
   41919: out<=1;
   41920: out<=1;
   41921: out<=0;
   41922: out<=0;
   41923: out<=1;
   41924: out<=0;
   41925: out<=0;
   41926: out<=0;
   41927: out<=0;
   41928: out<=0;
   41929: out<=0;
   41930: out<=1;
   41931: out<=1;
   41932: out<=1;
   41933: out<=0;
   41934: out<=1;
   41935: out<=0;
   41936: out<=0;
   41937: out<=0;
   41938: out<=0;
   41939: out<=0;
   41940: out<=0;
   41941: out<=1;
   41942: out<=1;
   41943: out<=0;
   41944: out<=0;
   41945: out<=1;
   41946: out<=0;
   41947: out<=1;
   41948: out<=0;
   41949: out<=0;
   41950: out<=1;
   41951: out<=1;
   41952: out<=1;
   41953: out<=1;
   41954: out<=0;
   41955: out<=0;
   41956: out<=1;
   41957: out<=0;
   41958: out<=1;
   41959: out<=0;
   41960: out<=0;
   41961: out<=1;
   41962: out<=1;
   41963: out<=0;
   41964: out<=0;
   41965: out<=0;
   41966: out<=0;
   41967: out<=0;
   41968: out<=0;
   41969: out<=1;
   41970: out<=0;
   41971: out<=1;
   41972: out<=1;
   41973: out<=1;
   41974: out<=0;
   41975: out<=0;
   41976: out<=0;
   41977: out<=0;
   41978: out<=0;
   41979: out<=0;
   41980: out<=1;
   41981: out<=0;
   41982: out<=0;
   41983: out<=1;
   41984: out<=0;
   41985: out<=0;
   41986: out<=1;
   41987: out<=1;
   41988: out<=1;
   41989: out<=0;
   41990: out<=1;
   41991: out<=0;
   41992: out<=0;
   41993: out<=1;
   41994: out<=1;
   41995: out<=0;
   41996: out<=1;
   41997: out<=1;
   41998: out<=1;
   41999: out<=1;
   42000: out<=1;
   42001: out<=0;
   42002: out<=1;
   42003: out<=0;
   42004: out<=1;
   42005: out<=1;
   42006: out<=0;
   42007: out<=0;
   42008: out<=0;
   42009: out<=0;
   42010: out<=0;
   42011: out<=0;
   42012: out<=0;
   42013: out<=1;
   42014: out<=1;
   42015: out<=0;
   42016: out<=0;
   42017: out<=1;
   42018: out<=1;
   42019: out<=0;
   42020: out<=0;
   42021: out<=0;
   42022: out<=0;
   42023: out<=0;
   42024: out<=0;
   42025: out<=0;
   42026: out<=1;
   42027: out<=1;
   42028: out<=0;
   42029: out<=1;
   42030: out<=0;
   42031: out<=1;
   42032: out<=1;
   42033: out<=1;
   42034: out<=1;
   42035: out<=1;
   42036: out<=0;
   42037: out<=1;
   42038: out<=1;
   42039: out<=0;
   42040: out<=0;
   42041: out<=1;
   42042: out<=0;
   42043: out<=1;
   42044: out<=1;
   42045: out<=1;
   42046: out<=0;
   42047: out<=0;
   42048: out<=1;
   42049: out<=1;
   42050: out<=0;
   42051: out<=0;
   42052: out<=0;
   42053: out<=1;
   42054: out<=0;
   42055: out<=1;
   42056: out<=1;
   42057: out<=0;
   42058: out<=0;
   42059: out<=1;
   42060: out<=0;
   42061: out<=0;
   42062: out<=0;
   42063: out<=0;
   42064: out<=1;
   42065: out<=0;
   42066: out<=1;
   42067: out<=0;
   42068: out<=1;
   42069: out<=1;
   42070: out<=0;
   42071: out<=0;
   42072: out<=0;
   42073: out<=0;
   42074: out<=0;
   42075: out<=0;
   42076: out<=0;
   42077: out<=1;
   42078: out<=1;
   42079: out<=0;
   42080: out<=0;
   42081: out<=1;
   42082: out<=1;
   42083: out<=0;
   42084: out<=0;
   42085: out<=0;
   42086: out<=0;
   42087: out<=0;
   42088: out<=0;
   42089: out<=0;
   42090: out<=1;
   42091: out<=1;
   42092: out<=0;
   42093: out<=1;
   42094: out<=0;
   42095: out<=1;
   42096: out<=0;
   42097: out<=0;
   42098: out<=0;
   42099: out<=0;
   42100: out<=1;
   42101: out<=0;
   42102: out<=0;
   42103: out<=1;
   42104: out<=1;
   42105: out<=0;
   42106: out<=1;
   42107: out<=0;
   42108: out<=0;
   42109: out<=0;
   42110: out<=1;
   42111: out<=1;
   42112: out<=1;
   42113: out<=1;
   42114: out<=0;
   42115: out<=0;
   42116: out<=0;
   42117: out<=1;
   42118: out<=0;
   42119: out<=1;
   42120: out<=1;
   42121: out<=0;
   42122: out<=0;
   42123: out<=1;
   42124: out<=0;
   42125: out<=0;
   42126: out<=0;
   42127: out<=0;
   42128: out<=1;
   42129: out<=0;
   42130: out<=1;
   42131: out<=0;
   42132: out<=1;
   42133: out<=1;
   42134: out<=0;
   42135: out<=0;
   42136: out<=0;
   42137: out<=0;
   42138: out<=0;
   42139: out<=0;
   42140: out<=0;
   42141: out<=1;
   42142: out<=1;
   42143: out<=0;
   42144: out<=1;
   42145: out<=0;
   42146: out<=0;
   42147: out<=1;
   42148: out<=1;
   42149: out<=1;
   42150: out<=1;
   42151: out<=1;
   42152: out<=1;
   42153: out<=1;
   42154: out<=0;
   42155: out<=0;
   42156: out<=1;
   42157: out<=0;
   42158: out<=1;
   42159: out<=0;
   42160: out<=1;
   42161: out<=1;
   42162: out<=1;
   42163: out<=1;
   42164: out<=0;
   42165: out<=1;
   42166: out<=1;
   42167: out<=0;
   42168: out<=0;
   42169: out<=1;
   42170: out<=0;
   42171: out<=1;
   42172: out<=1;
   42173: out<=1;
   42174: out<=0;
   42175: out<=0;
   42176: out<=0;
   42177: out<=0;
   42178: out<=1;
   42179: out<=1;
   42180: out<=1;
   42181: out<=0;
   42182: out<=1;
   42183: out<=0;
   42184: out<=0;
   42185: out<=1;
   42186: out<=1;
   42187: out<=0;
   42188: out<=1;
   42189: out<=1;
   42190: out<=1;
   42191: out<=1;
   42192: out<=1;
   42193: out<=0;
   42194: out<=1;
   42195: out<=0;
   42196: out<=1;
   42197: out<=1;
   42198: out<=0;
   42199: out<=0;
   42200: out<=0;
   42201: out<=0;
   42202: out<=0;
   42203: out<=0;
   42204: out<=0;
   42205: out<=1;
   42206: out<=1;
   42207: out<=0;
   42208: out<=1;
   42209: out<=0;
   42210: out<=0;
   42211: out<=1;
   42212: out<=1;
   42213: out<=1;
   42214: out<=1;
   42215: out<=1;
   42216: out<=1;
   42217: out<=1;
   42218: out<=0;
   42219: out<=0;
   42220: out<=1;
   42221: out<=0;
   42222: out<=1;
   42223: out<=0;
   42224: out<=0;
   42225: out<=0;
   42226: out<=0;
   42227: out<=0;
   42228: out<=1;
   42229: out<=0;
   42230: out<=0;
   42231: out<=1;
   42232: out<=1;
   42233: out<=0;
   42234: out<=1;
   42235: out<=0;
   42236: out<=0;
   42237: out<=0;
   42238: out<=1;
   42239: out<=1;
   42240: out<=1;
   42241: out<=0;
   42242: out<=1;
   42243: out<=0;
   42244: out<=1;
   42245: out<=1;
   42246: out<=0;
   42247: out<=0;
   42248: out<=0;
   42249: out<=0;
   42250: out<=0;
   42251: out<=0;
   42252: out<=0;
   42253: out<=1;
   42254: out<=1;
   42255: out<=0;
   42256: out<=1;
   42257: out<=1;
   42258: out<=0;
   42259: out<=0;
   42260: out<=0;
   42261: out<=1;
   42262: out<=0;
   42263: out<=1;
   42264: out<=1;
   42265: out<=0;
   42266: out<=0;
   42267: out<=1;
   42268: out<=0;
   42269: out<=0;
   42270: out<=0;
   42271: out<=0;
   42272: out<=0;
   42273: out<=0;
   42274: out<=0;
   42275: out<=0;
   42276: out<=1;
   42277: out<=0;
   42278: out<=0;
   42279: out<=1;
   42280: out<=1;
   42281: out<=0;
   42282: out<=1;
   42283: out<=0;
   42284: out<=0;
   42285: out<=0;
   42286: out<=1;
   42287: out<=1;
   42288: out<=0;
   42289: out<=1;
   42290: out<=1;
   42291: out<=0;
   42292: out<=0;
   42293: out<=0;
   42294: out<=0;
   42295: out<=0;
   42296: out<=0;
   42297: out<=0;
   42298: out<=1;
   42299: out<=1;
   42300: out<=0;
   42301: out<=1;
   42302: out<=0;
   42303: out<=1;
   42304: out<=1;
   42305: out<=0;
   42306: out<=1;
   42307: out<=0;
   42308: out<=1;
   42309: out<=1;
   42310: out<=0;
   42311: out<=0;
   42312: out<=0;
   42313: out<=0;
   42314: out<=0;
   42315: out<=0;
   42316: out<=0;
   42317: out<=1;
   42318: out<=1;
   42319: out<=0;
   42320: out<=0;
   42321: out<=0;
   42322: out<=1;
   42323: out<=1;
   42324: out<=1;
   42325: out<=0;
   42326: out<=1;
   42327: out<=0;
   42328: out<=0;
   42329: out<=1;
   42330: out<=1;
   42331: out<=0;
   42332: out<=1;
   42333: out<=1;
   42334: out<=1;
   42335: out<=1;
   42336: out<=1;
   42337: out<=1;
   42338: out<=1;
   42339: out<=1;
   42340: out<=0;
   42341: out<=1;
   42342: out<=1;
   42343: out<=0;
   42344: out<=0;
   42345: out<=1;
   42346: out<=0;
   42347: out<=1;
   42348: out<=1;
   42349: out<=1;
   42350: out<=0;
   42351: out<=0;
   42352: out<=0;
   42353: out<=1;
   42354: out<=1;
   42355: out<=0;
   42356: out<=0;
   42357: out<=0;
   42358: out<=0;
   42359: out<=0;
   42360: out<=0;
   42361: out<=0;
   42362: out<=1;
   42363: out<=1;
   42364: out<=0;
   42365: out<=1;
   42366: out<=0;
   42367: out<=1;
   42368: out<=1;
   42369: out<=0;
   42370: out<=1;
   42371: out<=0;
   42372: out<=1;
   42373: out<=1;
   42374: out<=0;
   42375: out<=0;
   42376: out<=0;
   42377: out<=0;
   42378: out<=0;
   42379: out<=0;
   42380: out<=0;
   42381: out<=1;
   42382: out<=1;
   42383: out<=0;
   42384: out<=0;
   42385: out<=0;
   42386: out<=1;
   42387: out<=1;
   42388: out<=1;
   42389: out<=0;
   42390: out<=1;
   42391: out<=0;
   42392: out<=0;
   42393: out<=1;
   42394: out<=1;
   42395: out<=0;
   42396: out<=1;
   42397: out<=1;
   42398: out<=1;
   42399: out<=1;
   42400: out<=0;
   42401: out<=0;
   42402: out<=0;
   42403: out<=0;
   42404: out<=1;
   42405: out<=0;
   42406: out<=0;
   42407: out<=1;
   42408: out<=1;
   42409: out<=0;
   42410: out<=1;
   42411: out<=0;
   42412: out<=0;
   42413: out<=0;
   42414: out<=1;
   42415: out<=1;
   42416: out<=1;
   42417: out<=0;
   42418: out<=0;
   42419: out<=1;
   42420: out<=1;
   42421: out<=1;
   42422: out<=1;
   42423: out<=1;
   42424: out<=1;
   42425: out<=1;
   42426: out<=0;
   42427: out<=0;
   42428: out<=1;
   42429: out<=0;
   42430: out<=1;
   42431: out<=0;
   42432: out<=1;
   42433: out<=0;
   42434: out<=1;
   42435: out<=0;
   42436: out<=1;
   42437: out<=1;
   42438: out<=0;
   42439: out<=0;
   42440: out<=0;
   42441: out<=0;
   42442: out<=0;
   42443: out<=0;
   42444: out<=0;
   42445: out<=1;
   42446: out<=1;
   42447: out<=0;
   42448: out<=1;
   42449: out<=1;
   42450: out<=0;
   42451: out<=0;
   42452: out<=0;
   42453: out<=1;
   42454: out<=0;
   42455: out<=1;
   42456: out<=1;
   42457: out<=0;
   42458: out<=0;
   42459: out<=1;
   42460: out<=0;
   42461: out<=0;
   42462: out<=0;
   42463: out<=0;
   42464: out<=1;
   42465: out<=1;
   42466: out<=1;
   42467: out<=1;
   42468: out<=0;
   42469: out<=1;
   42470: out<=1;
   42471: out<=0;
   42472: out<=0;
   42473: out<=1;
   42474: out<=0;
   42475: out<=1;
   42476: out<=1;
   42477: out<=1;
   42478: out<=0;
   42479: out<=0;
   42480: out<=1;
   42481: out<=0;
   42482: out<=0;
   42483: out<=1;
   42484: out<=1;
   42485: out<=1;
   42486: out<=1;
   42487: out<=1;
   42488: out<=1;
   42489: out<=1;
   42490: out<=0;
   42491: out<=0;
   42492: out<=1;
   42493: out<=0;
   42494: out<=1;
   42495: out<=0;
   42496: out<=1;
   42497: out<=0;
   42498: out<=0;
   42499: out<=1;
   42500: out<=1;
   42501: out<=1;
   42502: out<=1;
   42503: out<=1;
   42504: out<=1;
   42505: out<=1;
   42506: out<=0;
   42507: out<=0;
   42508: out<=1;
   42509: out<=0;
   42510: out<=1;
   42511: out<=0;
   42512: out<=1;
   42513: out<=1;
   42514: out<=1;
   42515: out<=1;
   42516: out<=0;
   42517: out<=1;
   42518: out<=1;
   42519: out<=0;
   42520: out<=0;
   42521: out<=1;
   42522: out<=0;
   42523: out<=1;
   42524: out<=1;
   42525: out<=1;
   42526: out<=0;
   42527: out<=0;
   42528: out<=1;
   42529: out<=1;
   42530: out<=0;
   42531: out<=0;
   42532: out<=0;
   42533: out<=1;
   42534: out<=0;
   42535: out<=1;
   42536: out<=1;
   42537: out<=0;
   42538: out<=0;
   42539: out<=1;
   42540: out<=0;
   42541: out<=0;
   42542: out<=0;
   42543: out<=0;
   42544: out<=1;
   42545: out<=0;
   42546: out<=1;
   42547: out<=0;
   42548: out<=1;
   42549: out<=1;
   42550: out<=0;
   42551: out<=0;
   42552: out<=0;
   42553: out<=0;
   42554: out<=0;
   42555: out<=0;
   42556: out<=0;
   42557: out<=1;
   42558: out<=1;
   42559: out<=0;
   42560: out<=1;
   42561: out<=0;
   42562: out<=0;
   42563: out<=1;
   42564: out<=1;
   42565: out<=1;
   42566: out<=1;
   42567: out<=1;
   42568: out<=1;
   42569: out<=1;
   42570: out<=0;
   42571: out<=0;
   42572: out<=1;
   42573: out<=0;
   42574: out<=1;
   42575: out<=0;
   42576: out<=0;
   42577: out<=0;
   42578: out<=0;
   42579: out<=0;
   42580: out<=1;
   42581: out<=0;
   42582: out<=0;
   42583: out<=1;
   42584: out<=1;
   42585: out<=0;
   42586: out<=1;
   42587: out<=0;
   42588: out<=0;
   42589: out<=0;
   42590: out<=1;
   42591: out<=1;
   42592: out<=0;
   42593: out<=0;
   42594: out<=1;
   42595: out<=1;
   42596: out<=1;
   42597: out<=0;
   42598: out<=1;
   42599: out<=0;
   42600: out<=0;
   42601: out<=1;
   42602: out<=1;
   42603: out<=0;
   42604: out<=1;
   42605: out<=1;
   42606: out<=1;
   42607: out<=1;
   42608: out<=1;
   42609: out<=0;
   42610: out<=1;
   42611: out<=0;
   42612: out<=1;
   42613: out<=1;
   42614: out<=0;
   42615: out<=0;
   42616: out<=0;
   42617: out<=0;
   42618: out<=0;
   42619: out<=0;
   42620: out<=0;
   42621: out<=1;
   42622: out<=1;
   42623: out<=0;
   42624: out<=0;
   42625: out<=1;
   42626: out<=1;
   42627: out<=0;
   42628: out<=0;
   42629: out<=0;
   42630: out<=0;
   42631: out<=0;
   42632: out<=0;
   42633: out<=0;
   42634: out<=1;
   42635: out<=1;
   42636: out<=0;
   42637: out<=1;
   42638: out<=0;
   42639: out<=1;
   42640: out<=1;
   42641: out<=1;
   42642: out<=1;
   42643: out<=1;
   42644: out<=0;
   42645: out<=1;
   42646: out<=1;
   42647: out<=0;
   42648: out<=0;
   42649: out<=1;
   42650: out<=0;
   42651: out<=1;
   42652: out<=1;
   42653: out<=1;
   42654: out<=0;
   42655: out<=0;
   42656: out<=0;
   42657: out<=0;
   42658: out<=1;
   42659: out<=1;
   42660: out<=1;
   42661: out<=0;
   42662: out<=1;
   42663: out<=0;
   42664: out<=0;
   42665: out<=1;
   42666: out<=1;
   42667: out<=0;
   42668: out<=1;
   42669: out<=1;
   42670: out<=1;
   42671: out<=1;
   42672: out<=1;
   42673: out<=0;
   42674: out<=1;
   42675: out<=0;
   42676: out<=1;
   42677: out<=1;
   42678: out<=0;
   42679: out<=0;
   42680: out<=0;
   42681: out<=0;
   42682: out<=0;
   42683: out<=0;
   42684: out<=0;
   42685: out<=1;
   42686: out<=1;
   42687: out<=0;
   42688: out<=0;
   42689: out<=1;
   42690: out<=1;
   42691: out<=0;
   42692: out<=0;
   42693: out<=0;
   42694: out<=0;
   42695: out<=0;
   42696: out<=0;
   42697: out<=0;
   42698: out<=1;
   42699: out<=1;
   42700: out<=0;
   42701: out<=1;
   42702: out<=0;
   42703: out<=1;
   42704: out<=0;
   42705: out<=0;
   42706: out<=0;
   42707: out<=0;
   42708: out<=1;
   42709: out<=0;
   42710: out<=0;
   42711: out<=1;
   42712: out<=1;
   42713: out<=0;
   42714: out<=1;
   42715: out<=0;
   42716: out<=0;
   42717: out<=0;
   42718: out<=1;
   42719: out<=1;
   42720: out<=1;
   42721: out<=1;
   42722: out<=0;
   42723: out<=0;
   42724: out<=0;
   42725: out<=1;
   42726: out<=0;
   42727: out<=1;
   42728: out<=1;
   42729: out<=0;
   42730: out<=0;
   42731: out<=1;
   42732: out<=0;
   42733: out<=0;
   42734: out<=0;
   42735: out<=0;
   42736: out<=1;
   42737: out<=0;
   42738: out<=1;
   42739: out<=0;
   42740: out<=1;
   42741: out<=1;
   42742: out<=0;
   42743: out<=0;
   42744: out<=0;
   42745: out<=0;
   42746: out<=0;
   42747: out<=0;
   42748: out<=0;
   42749: out<=1;
   42750: out<=1;
   42751: out<=0;
   42752: out<=0;
   42753: out<=0;
   42754: out<=0;
   42755: out<=0;
   42756: out<=1;
   42757: out<=0;
   42758: out<=0;
   42759: out<=1;
   42760: out<=1;
   42761: out<=0;
   42762: out<=1;
   42763: out<=0;
   42764: out<=0;
   42765: out<=0;
   42766: out<=1;
   42767: out<=1;
   42768: out<=1;
   42769: out<=0;
   42770: out<=0;
   42771: out<=1;
   42772: out<=1;
   42773: out<=1;
   42774: out<=1;
   42775: out<=1;
   42776: out<=1;
   42777: out<=1;
   42778: out<=0;
   42779: out<=0;
   42780: out<=1;
   42781: out<=0;
   42782: out<=1;
   42783: out<=0;
   42784: out<=1;
   42785: out<=0;
   42786: out<=1;
   42787: out<=0;
   42788: out<=1;
   42789: out<=1;
   42790: out<=0;
   42791: out<=0;
   42792: out<=0;
   42793: out<=0;
   42794: out<=0;
   42795: out<=0;
   42796: out<=0;
   42797: out<=1;
   42798: out<=1;
   42799: out<=0;
   42800: out<=0;
   42801: out<=0;
   42802: out<=1;
   42803: out<=1;
   42804: out<=1;
   42805: out<=0;
   42806: out<=1;
   42807: out<=0;
   42808: out<=0;
   42809: out<=1;
   42810: out<=1;
   42811: out<=0;
   42812: out<=1;
   42813: out<=1;
   42814: out<=1;
   42815: out<=1;
   42816: out<=1;
   42817: out<=1;
   42818: out<=1;
   42819: out<=1;
   42820: out<=0;
   42821: out<=1;
   42822: out<=1;
   42823: out<=0;
   42824: out<=0;
   42825: out<=1;
   42826: out<=0;
   42827: out<=1;
   42828: out<=1;
   42829: out<=1;
   42830: out<=0;
   42831: out<=0;
   42832: out<=1;
   42833: out<=0;
   42834: out<=0;
   42835: out<=1;
   42836: out<=1;
   42837: out<=1;
   42838: out<=1;
   42839: out<=1;
   42840: out<=1;
   42841: out<=1;
   42842: out<=0;
   42843: out<=0;
   42844: out<=1;
   42845: out<=0;
   42846: out<=1;
   42847: out<=0;
   42848: out<=1;
   42849: out<=0;
   42850: out<=1;
   42851: out<=0;
   42852: out<=1;
   42853: out<=1;
   42854: out<=0;
   42855: out<=0;
   42856: out<=0;
   42857: out<=0;
   42858: out<=0;
   42859: out<=0;
   42860: out<=0;
   42861: out<=1;
   42862: out<=1;
   42863: out<=0;
   42864: out<=1;
   42865: out<=1;
   42866: out<=0;
   42867: out<=0;
   42868: out<=0;
   42869: out<=1;
   42870: out<=0;
   42871: out<=1;
   42872: out<=1;
   42873: out<=0;
   42874: out<=0;
   42875: out<=1;
   42876: out<=0;
   42877: out<=0;
   42878: out<=0;
   42879: out<=0;
   42880: out<=0;
   42881: out<=0;
   42882: out<=0;
   42883: out<=0;
   42884: out<=1;
   42885: out<=0;
   42886: out<=0;
   42887: out<=1;
   42888: out<=1;
   42889: out<=0;
   42890: out<=1;
   42891: out<=0;
   42892: out<=0;
   42893: out<=0;
   42894: out<=1;
   42895: out<=1;
   42896: out<=0;
   42897: out<=1;
   42898: out<=1;
   42899: out<=0;
   42900: out<=0;
   42901: out<=0;
   42902: out<=0;
   42903: out<=0;
   42904: out<=0;
   42905: out<=0;
   42906: out<=1;
   42907: out<=1;
   42908: out<=0;
   42909: out<=1;
   42910: out<=0;
   42911: out<=1;
   42912: out<=1;
   42913: out<=0;
   42914: out<=1;
   42915: out<=0;
   42916: out<=1;
   42917: out<=1;
   42918: out<=0;
   42919: out<=0;
   42920: out<=0;
   42921: out<=0;
   42922: out<=0;
   42923: out<=0;
   42924: out<=0;
   42925: out<=1;
   42926: out<=1;
   42927: out<=0;
   42928: out<=1;
   42929: out<=1;
   42930: out<=0;
   42931: out<=0;
   42932: out<=0;
   42933: out<=1;
   42934: out<=0;
   42935: out<=1;
   42936: out<=1;
   42937: out<=0;
   42938: out<=0;
   42939: out<=1;
   42940: out<=0;
   42941: out<=0;
   42942: out<=0;
   42943: out<=0;
   42944: out<=1;
   42945: out<=1;
   42946: out<=1;
   42947: out<=1;
   42948: out<=0;
   42949: out<=1;
   42950: out<=1;
   42951: out<=0;
   42952: out<=0;
   42953: out<=1;
   42954: out<=0;
   42955: out<=1;
   42956: out<=1;
   42957: out<=1;
   42958: out<=0;
   42959: out<=0;
   42960: out<=0;
   42961: out<=1;
   42962: out<=1;
   42963: out<=0;
   42964: out<=0;
   42965: out<=0;
   42966: out<=0;
   42967: out<=0;
   42968: out<=0;
   42969: out<=0;
   42970: out<=1;
   42971: out<=1;
   42972: out<=0;
   42973: out<=1;
   42974: out<=0;
   42975: out<=1;
   42976: out<=1;
   42977: out<=0;
   42978: out<=1;
   42979: out<=0;
   42980: out<=1;
   42981: out<=1;
   42982: out<=0;
   42983: out<=0;
   42984: out<=0;
   42985: out<=0;
   42986: out<=0;
   42987: out<=0;
   42988: out<=0;
   42989: out<=1;
   42990: out<=1;
   42991: out<=0;
   42992: out<=0;
   42993: out<=0;
   42994: out<=1;
   42995: out<=1;
   42996: out<=1;
   42997: out<=0;
   42998: out<=1;
   42999: out<=0;
   43000: out<=0;
   43001: out<=1;
   43002: out<=1;
   43003: out<=0;
   43004: out<=1;
   43005: out<=1;
   43006: out<=1;
   43007: out<=1;
   43008: out<=0;
   43009: out<=0;
   43010: out<=0;
   43011: out<=0;
   43012: out<=1;
   43013: out<=0;
   43014: out<=0;
   43015: out<=1;
   43016: out<=0;
   43017: out<=1;
   43018: out<=0;
   43019: out<=1;
   43020: out<=1;
   43021: out<=1;
   43022: out<=0;
   43023: out<=0;
   43024: out<=1;
   43025: out<=0;
   43026: out<=0;
   43027: out<=1;
   43028: out<=1;
   43029: out<=1;
   43030: out<=1;
   43031: out<=1;
   43032: out<=0;
   43033: out<=0;
   43034: out<=1;
   43035: out<=1;
   43036: out<=0;
   43037: out<=1;
   43038: out<=0;
   43039: out<=1;
   43040: out<=0;
   43041: out<=1;
   43042: out<=0;
   43043: out<=1;
   43044: out<=0;
   43045: out<=0;
   43046: out<=1;
   43047: out<=1;
   43048: out<=0;
   43049: out<=0;
   43050: out<=0;
   43051: out<=0;
   43052: out<=0;
   43053: out<=1;
   43054: out<=1;
   43055: out<=0;
   43056: out<=1;
   43057: out<=1;
   43058: out<=0;
   43059: out<=0;
   43060: out<=0;
   43061: out<=1;
   43062: out<=0;
   43063: out<=1;
   43064: out<=0;
   43065: out<=1;
   43066: out<=1;
   43067: out<=0;
   43068: out<=1;
   43069: out<=1;
   43070: out<=1;
   43071: out<=1;
   43072: out<=1;
   43073: out<=1;
   43074: out<=1;
   43075: out<=1;
   43076: out<=0;
   43077: out<=1;
   43078: out<=1;
   43079: out<=0;
   43080: out<=1;
   43081: out<=0;
   43082: out<=1;
   43083: out<=0;
   43084: out<=0;
   43085: out<=0;
   43086: out<=1;
   43087: out<=1;
   43088: out<=1;
   43089: out<=0;
   43090: out<=0;
   43091: out<=1;
   43092: out<=1;
   43093: out<=1;
   43094: out<=1;
   43095: out<=1;
   43096: out<=0;
   43097: out<=0;
   43098: out<=1;
   43099: out<=1;
   43100: out<=0;
   43101: out<=1;
   43102: out<=0;
   43103: out<=1;
   43104: out<=0;
   43105: out<=1;
   43106: out<=0;
   43107: out<=1;
   43108: out<=0;
   43109: out<=0;
   43110: out<=1;
   43111: out<=1;
   43112: out<=0;
   43113: out<=0;
   43114: out<=0;
   43115: out<=0;
   43116: out<=0;
   43117: out<=1;
   43118: out<=1;
   43119: out<=0;
   43120: out<=0;
   43121: out<=0;
   43122: out<=1;
   43123: out<=1;
   43124: out<=1;
   43125: out<=0;
   43126: out<=1;
   43127: out<=0;
   43128: out<=1;
   43129: out<=0;
   43130: out<=0;
   43131: out<=1;
   43132: out<=0;
   43133: out<=0;
   43134: out<=0;
   43135: out<=0;
   43136: out<=0;
   43137: out<=0;
   43138: out<=0;
   43139: out<=0;
   43140: out<=1;
   43141: out<=0;
   43142: out<=0;
   43143: out<=1;
   43144: out<=0;
   43145: out<=1;
   43146: out<=0;
   43147: out<=1;
   43148: out<=1;
   43149: out<=1;
   43150: out<=0;
   43151: out<=0;
   43152: out<=0;
   43153: out<=1;
   43154: out<=1;
   43155: out<=0;
   43156: out<=0;
   43157: out<=0;
   43158: out<=0;
   43159: out<=0;
   43160: out<=1;
   43161: out<=1;
   43162: out<=0;
   43163: out<=0;
   43164: out<=1;
   43165: out<=0;
   43166: out<=1;
   43167: out<=0;
   43168: out<=0;
   43169: out<=1;
   43170: out<=0;
   43171: out<=1;
   43172: out<=0;
   43173: out<=0;
   43174: out<=1;
   43175: out<=1;
   43176: out<=0;
   43177: out<=0;
   43178: out<=0;
   43179: out<=0;
   43180: out<=0;
   43181: out<=1;
   43182: out<=1;
   43183: out<=0;
   43184: out<=0;
   43185: out<=0;
   43186: out<=1;
   43187: out<=1;
   43188: out<=1;
   43189: out<=0;
   43190: out<=1;
   43191: out<=0;
   43192: out<=1;
   43193: out<=0;
   43194: out<=0;
   43195: out<=1;
   43196: out<=0;
   43197: out<=0;
   43198: out<=0;
   43199: out<=0;
   43200: out<=1;
   43201: out<=1;
   43202: out<=1;
   43203: out<=1;
   43204: out<=0;
   43205: out<=1;
   43206: out<=1;
   43207: out<=0;
   43208: out<=1;
   43209: out<=0;
   43210: out<=1;
   43211: out<=0;
   43212: out<=0;
   43213: out<=0;
   43214: out<=1;
   43215: out<=1;
   43216: out<=0;
   43217: out<=1;
   43218: out<=1;
   43219: out<=0;
   43220: out<=0;
   43221: out<=0;
   43222: out<=0;
   43223: out<=0;
   43224: out<=1;
   43225: out<=1;
   43226: out<=0;
   43227: out<=0;
   43228: out<=1;
   43229: out<=0;
   43230: out<=1;
   43231: out<=0;
   43232: out<=0;
   43233: out<=1;
   43234: out<=0;
   43235: out<=1;
   43236: out<=0;
   43237: out<=0;
   43238: out<=1;
   43239: out<=1;
   43240: out<=0;
   43241: out<=0;
   43242: out<=0;
   43243: out<=0;
   43244: out<=0;
   43245: out<=1;
   43246: out<=1;
   43247: out<=0;
   43248: out<=1;
   43249: out<=1;
   43250: out<=0;
   43251: out<=0;
   43252: out<=0;
   43253: out<=1;
   43254: out<=0;
   43255: out<=1;
   43256: out<=0;
   43257: out<=1;
   43258: out<=1;
   43259: out<=0;
   43260: out<=1;
   43261: out<=1;
   43262: out<=1;
   43263: out<=1;
   43264: out<=1;
   43265: out<=0;
   43266: out<=0;
   43267: out<=1;
   43268: out<=1;
   43269: out<=1;
   43270: out<=1;
   43271: out<=1;
   43272: out<=0;
   43273: out<=0;
   43274: out<=1;
   43275: out<=1;
   43276: out<=0;
   43277: out<=1;
   43278: out<=0;
   43279: out<=1;
   43280: out<=1;
   43281: out<=1;
   43282: out<=1;
   43283: out<=1;
   43284: out<=0;
   43285: out<=1;
   43286: out<=1;
   43287: out<=0;
   43288: out<=1;
   43289: out<=0;
   43290: out<=1;
   43291: out<=0;
   43292: out<=0;
   43293: out<=0;
   43294: out<=1;
   43295: out<=1;
   43296: out<=0;
   43297: out<=0;
   43298: out<=1;
   43299: out<=1;
   43300: out<=1;
   43301: out<=0;
   43302: out<=1;
   43303: out<=0;
   43304: out<=1;
   43305: out<=0;
   43306: out<=0;
   43307: out<=1;
   43308: out<=0;
   43309: out<=0;
   43310: out<=0;
   43311: out<=0;
   43312: out<=0;
   43313: out<=1;
   43314: out<=0;
   43315: out<=1;
   43316: out<=0;
   43317: out<=0;
   43318: out<=1;
   43319: out<=1;
   43320: out<=0;
   43321: out<=0;
   43322: out<=0;
   43323: out<=0;
   43324: out<=0;
   43325: out<=1;
   43326: out<=1;
   43327: out<=0;
   43328: out<=1;
   43329: out<=0;
   43330: out<=0;
   43331: out<=1;
   43332: out<=1;
   43333: out<=1;
   43334: out<=1;
   43335: out<=1;
   43336: out<=0;
   43337: out<=0;
   43338: out<=1;
   43339: out<=1;
   43340: out<=0;
   43341: out<=1;
   43342: out<=0;
   43343: out<=1;
   43344: out<=0;
   43345: out<=0;
   43346: out<=0;
   43347: out<=0;
   43348: out<=1;
   43349: out<=0;
   43350: out<=0;
   43351: out<=1;
   43352: out<=0;
   43353: out<=1;
   43354: out<=0;
   43355: out<=1;
   43356: out<=1;
   43357: out<=1;
   43358: out<=0;
   43359: out<=0;
   43360: out<=1;
   43361: out<=1;
   43362: out<=0;
   43363: out<=0;
   43364: out<=0;
   43365: out<=1;
   43366: out<=0;
   43367: out<=1;
   43368: out<=0;
   43369: out<=1;
   43370: out<=1;
   43371: out<=0;
   43372: out<=1;
   43373: out<=1;
   43374: out<=1;
   43375: out<=1;
   43376: out<=0;
   43377: out<=1;
   43378: out<=0;
   43379: out<=1;
   43380: out<=0;
   43381: out<=0;
   43382: out<=1;
   43383: out<=1;
   43384: out<=0;
   43385: out<=0;
   43386: out<=0;
   43387: out<=0;
   43388: out<=0;
   43389: out<=1;
   43390: out<=1;
   43391: out<=0;
   43392: out<=0;
   43393: out<=1;
   43394: out<=1;
   43395: out<=0;
   43396: out<=0;
   43397: out<=0;
   43398: out<=0;
   43399: out<=0;
   43400: out<=1;
   43401: out<=1;
   43402: out<=0;
   43403: out<=0;
   43404: out<=1;
   43405: out<=0;
   43406: out<=1;
   43407: out<=0;
   43408: out<=1;
   43409: out<=1;
   43410: out<=1;
   43411: out<=1;
   43412: out<=0;
   43413: out<=1;
   43414: out<=1;
   43415: out<=0;
   43416: out<=1;
   43417: out<=0;
   43418: out<=1;
   43419: out<=0;
   43420: out<=0;
   43421: out<=0;
   43422: out<=1;
   43423: out<=1;
   43424: out<=1;
   43425: out<=1;
   43426: out<=0;
   43427: out<=0;
   43428: out<=0;
   43429: out<=1;
   43430: out<=0;
   43431: out<=1;
   43432: out<=0;
   43433: out<=1;
   43434: out<=1;
   43435: out<=0;
   43436: out<=1;
   43437: out<=1;
   43438: out<=1;
   43439: out<=1;
   43440: out<=0;
   43441: out<=1;
   43442: out<=0;
   43443: out<=1;
   43444: out<=0;
   43445: out<=0;
   43446: out<=1;
   43447: out<=1;
   43448: out<=0;
   43449: out<=0;
   43450: out<=0;
   43451: out<=0;
   43452: out<=0;
   43453: out<=1;
   43454: out<=1;
   43455: out<=0;
   43456: out<=0;
   43457: out<=1;
   43458: out<=1;
   43459: out<=0;
   43460: out<=0;
   43461: out<=0;
   43462: out<=0;
   43463: out<=0;
   43464: out<=1;
   43465: out<=1;
   43466: out<=0;
   43467: out<=0;
   43468: out<=1;
   43469: out<=0;
   43470: out<=1;
   43471: out<=0;
   43472: out<=0;
   43473: out<=0;
   43474: out<=0;
   43475: out<=0;
   43476: out<=1;
   43477: out<=0;
   43478: out<=0;
   43479: out<=1;
   43480: out<=0;
   43481: out<=1;
   43482: out<=0;
   43483: out<=1;
   43484: out<=1;
   43485: out<=1;
   43486: out<=0;
   43487: out<=0;
   43488: out<=0;
   43489: out<=0;
   43490: out<=1;
   43491: out<=1;
   43492: out<=1;
   43493: out<=0;
   43494: out<=1;
   43495: out<=0;
   43496: out<=1;
   43497: out<=0;
   43498: out<=0;
   43499: out<=1;
   43500: out<=0;
   43501: out<=0;
   43502: out<=0;
   43503: out<=0;
   43504: out<=0;
   43505: out<=1;
   43506: out<=0;
   43507: out<=1;
   43508: out<=0;
   43509: out<=0;
   43510: out<=1;
   43511: out<=1;
   43512: out<=0;
   43513: out<=0;
   43514: out<=0;
   43515: out<=0;
   43516: out<=0;
   43517: out<=1;
   43518: out<=1;
   43519: out<=0;
   43520: out<=0;
   43521: out<=1;
   43522: out<=0;
   43523: out<=1;
   43524: out<=0;
   43525: out<=0;
   43526: out<=1;
   43527: out<=1;
   43528: out<=0;
   43529: out<=0;
   43530: out<=0;
   43531: out<=0;
   43532: out<=0;
   43533: out<=1;
   43534: out<=1;
   43535: out<=0;
   43536: out<=0;
   43537: out<=0;
   43538: out<=1;
   43539: out<=1;
   43540: out<=1;
   43541: out<=0;
   43542: out<=1;
   43543: out<=0;
   43544: out<=1;
   43545: out<=0;
   43546: out<=0;
   43547: out<=1;
   43548: out<=0;
   43549: out<=0;
   43550: out<=0;
   43551: out<=0;
   43552: out<=0;
   43553: out<=0;
   43554: out<=0;
   43555: out<=0;
   43556: out<=1;
   43557: out<=0;
   43558: out<=0;
   43559: out<=1;
   43560: out<=0;
   43561: out<=1;
   43562: out<=0;
   43563: out<=1;
   43564: out<=1;
   43565: out<=1;
   43566: out<=0;
   43567: out<=0;
   43568: out<=0;
   43569: out<=1;
   43570: out<=1;
   43571: out<=0;
   43572: out<=0;
   43573: out<=0;
   43574: out<=0;
   43575: out<=0;
   43576: out<=1;
   43577: out<=1;
   43578: out<=0;
   43579: out<=0;
   43580: out<=1;
   43581: out<=0;
   43582: out<=1;
   43583: out<=0;
   43584: out<=0;
   43585: out<=1;
   43586: out<=0;
   43587: out<=1;
   43588: out<=0;
   43589: out<=0;
   43590: out<=1;
   43591: out<=1;
   43592: out<=0;
   43593: out<=0;
   43594: out<=0;
   43595: out<=0;
   43596: out<=0;
   43597: out<=1;
   43598: out<=1;
   43599: out<=0;
   43600: out<=1;
   43601: out<=1;
   43602: out<=0;
   43603: out<=0;
   43604: out<=0;
   43605: out<=1;
   43606: out<=0;
   43607: out<=1;
   43608: out<=0;
   43609: out<=1;
   43610: out<=1;
   43611: out<=0;
   43612: out<=1;
   43613: out<=1;
   43614: out<=1;
   43615: out<=1;
   43616: out<=1;
   43617: out<=1;
   43618: out<=1;
   43619: out<=1;
   43620: out<=0;
   43621: out<=1;
   43622: out<=1;
   43623: out<=0;
   43624: out<=1;
   43625: out<=0;
   43626: out<=1;
   43627: out<=0;
   43628: out<=0;
   43629: out<=0;
   43630: out<=1;
   43631: out<=1;
   43632: out<=0;
   43633: out<=1;
   43634: out<=1;
   43635: out<=0;
   43636: out<=0;
   43637: out<=0;
   43638: out<=0;
   43639: out<=0;
   43640: out<=1;
   43641: out<=1;
   43642: out<=0;
   43643: out<=0;
   43644: out<=1;
   43645: out<=0;
   43646: out<=1;
   43647: out<=0;
   43648: out<=0;
   43649: out<=1;
   43650: out<=0;
   43651: out<=1;
   43652: out<=0;
   43653: out<=0;
   43654: out<=1;
   43655: out<=1;
   43656: out<=0;
   43657: out<=0;
   43658: out<=0;
   43659: out<=0;
   43660: out<=0;
   43661: out<=1;
   43662: out<=1;
   43663: out<=0;
   43664: out<=1;
   43665: out<=1;
   43666: out<=0;
   43667: out<=0;
   43668: out<=0;
   43669: out<=1;
   43670: out<=0;
   43671: out<=1;
   43672: out<=0;
   43673: out<=1;
   43674: out<=1;
   43675: out<=0;
   43676: out<=1;
   43677: out<=1;
   43678: out<=1;
   43679: out<=1;
   43680: out<=0;
   43681: out<=0;
   43682: out<=0;
   43683: out<=0;
   43684: out<=1;
   43685: out<=0;
   43686: out<=0;
   43687: out<=1;
   43688: out<=0;
   43689: out<=1;
   43690: out<=0;
   43691: out<=1;
   43692: out<=1;
   43693: out<=1;
   43694: out<=0;
   43695: out<=0;
   43696: out<=1;
   43697: out<=0;
   43698: out<=0;
   43699: out<=1;
   43700: out<=1;
   43701: out<=1;
   43702: out<=1;
   43703: out<=1;
   43704: out<=0;
   43705: out<=0;
   43706: out<=1;
   43707: out<=1;
   43708: out<=0;
   43709: out<=1;
   43710: out<=0;
   43711: out<=1;
   43712: out<=0;
   43713: out<=1;
   43714: out<=0;
   43715: out<=1;
   43716: out<=0;
   43717: out<=0;
   43718: out<=1;
   43719: out<=1;
   43720: out<=0;
   43721: out<=0;
   43722: out<=0;
   43723: out<=0;
   43724: out<=0;
   43725: out<=1;
   43726: out<=1;
   43727: out<=0;
   43728: out<=0;
   43729: out<=0;
   43730: out<=1;
   43731: out<=1;
   43732: out<=1;
   43733: out<=0;
   43734: out<=1;
   43735: out<=0;
   43736: out<=1;
   43737: out<=0;
   43738: out<=0;
   43739: out<=1;
   43740: out<=0;
   43741: out<=0;
   43742: out<=0;
   43743: out<=0;
   43744: out<=1;
   43745: out<=1;
   43746: out<=1;
   43747: out<=1;
   43748: out<=0;
   43749: out<=1;
   43750: out<=1;
   43751: out<=0;
   43752: out<=1;
   43753: out<=0;
   43754: out<=1;
   43755: out<=0;
   43756: out<=0;
   43757: out<=0;
   43758: out<=1;
   43759: out<=1;
   43760: out<=1;
   43761: out<=0;
   43762: out<=0;
   43763: out<=1;
   43764: out<=1;
   43765: out<=1;
   43766: out<=1;
   43767: out<=1;
   43768: out<=0;
   43769: out<=0;
   43770: out<=1;
   43771: out<=1;
   43772: out<=0;
   43773: out<=1;
   43774: out<=0;
   43775: out<=1;
   43776: out<=1;
   43777: out<=1;
   43778: out<=0;
   43779: out<=0;
   43780: out<=0;
   43781: out<=1;
   43782: out<=0;
   43783: out<=1;
   43784: out<=0;
   43785: out<=1;
   43786: out<=1;
   43787: out<=0;
   43788: out<=1;
   43789: out<=1;
   43790: out<=1;
   43791: out<=1;
   43792: out<=0;
   43793: out<=1;
   43794: out<=0;
   43795: out<=1;
   43796: out<=0;
   43797: out<=0;
   43798: out<=1;
   43799: out<=1;
   43800: out<=0;
   43801: out<=0;
   43802: out<=0;
   43803: out<=0;
   43804: out<=0;
   43805: out<=1;
   43806: out<=1;
   43807: out<=0;
   43808: out<=0;
   43809: out<=1;
   43810: out<=1;
   43811: out<=0;
   43812: out<=0;
   43813: out<=0;
   43814: out<=0;
   43815: out<=0;
   43816: out<=1;
   43817: out<=1;
   43818: out<=0;
   43819: out<=0;
   43820: out<=1;
   43821: out<=0;
   43822: out<=1;
   43823: out<=0;
   43824: out<=1;
   43825: out<=1;
   43826: out<=1;
   43827: out<=1;
   43828: out<=0;
   43829: out<=1;
   43830: out<=1;
   43831: out<=0;
   43832: out<=1;
   43833: out<=0;
   43834: out<=1;
   43835: out<=0;
   43836: out<=0;
   43837: out<=0;
   43838: out<=1;
   43839: out<=1;
   43840: out<=0;
   43841: out<=0;
   43842: out<=1;
   43843: out<=1;
   43844: out<=1;
   43845: out<=0;
   43846: out<=1;
   43847: out<=0;
   43848: out<=1;
   43849: out<=0;
   43850: out<=0;
   43851: out<=1;
   43852: out<=0;
   43853: out<=0;
   43854: out<=0;
   43855: out<=0;
   43856: out<=0;
   43857: out<=1;
   43858: out<=0;
   43859: out<=1;
   43860: out<=0;
   43861: out<=0;
   43862: out<=1;
   43863: out<=1;
   43864: out<=0;
   43865: out<=0;
   43866: out<=0;
   43867: out<=0;
   43868: out<=0;
   43869: out<=1;
   43870: out<=1;
   43871: out<=0;
   43872: out<=0;
   43873: out<=1;
   43874: out<=1;
   43875: out<=0;
   43876: out<=0;
   43877: out<=0;
   43878: out<=0;
   43879: out<=0;
   43880: out<=1;
   43881: out<=1;
   43882: out<=0;
   43883: out<=0;
   43884: out<=1;
   43885: out<=0;
   43886: out<=1;
   43887: out<=0;
   43888: out<=0;
   43889: out<=0;
   43890: out<=0;
   43891: out<=0;
   43892: out<=1;
   43893: out<=0;
   43894: out<=0;
   43895: out<=1;
   43896: out<=0;
   43897: out<=1;
   43898: out<=0;
   43899: out<=1;
   43900: out<=1;
   43901: out<=1;
   43902: out<=0;
   43903: out<=0;
   43904: out<=0;
   43905: out<=0;
   43906: out<=1;
   43907: out<=1;
   43908: out<=1;
   43909: out<=0;
   43910: out<=1;
   43911: out<=0;
   43912: out<=1;
   43913: out<=0;
   43914: out<=0;
   43915: out<=1;
   43916: out<=0;
   43917: out<=0;
   43918: out<=0;
   43919: out<=0;
   43920: out<=0;
   43921: out<=1;
   43922: out<=0;
   43923: out<=1;
   43924: out<=0;
   43925: out<=0;
   43926: out<=1;
   43927: out<=1;
   43928: out<=0;
   43929: out<=0;
   43930: out<=0;
   43931: out<=0;
   43932: out<=0;
   43933: out<=1;
   43934: out<=1;
   43935: out<=0;
   43936: out<=1;
   43937: out<=0;
   43938: out<=0;
   43939: out<=1;
   43940: out<=1;
   43941: out<=1;
   43942: out<=1;
   43943: out<=1;
   43944: out<=0;
   43945: out<=0;
   43946: out<=1;
   43947: out<=1;
   43948: out<=0;
   43949: out<=1;
   43950: out<=0;
   43951: out<=1;
   43952: out<=1;
   43953: out<=1;
   43954: out<=1;
   43955: out<=1;
   43956: out<=0;
   43957: out<=1;
   43958: out<=1;
   43959: out<=0;
   43960: out<=1;
   43961: out<=0;
   43962: out<=1;
   43963: out<=0;
   43964: out<=0;
   43965: out<=0;
   43966: out<=1;
   43967: out<=1;
   43968: out<=1;
   43969: out<=1;
   43970: out<=0;
   43971: out<=0;
   43972: out<=0;
   43973: out<=1;
   43974: out<=0;
   43975: out<=1;
   43976: out<=0;
   43977: out<=1;
   43978: out<=1;
   43979: out<=0;
   43980: out<=1;
   43981: out<=1;
   43982: out<=1;
   43983: out<=1;
   43984: out<=0;
   43985: out<=1;
   43986: out<=0;
   43987: out<=1;
   43988: out<=0;
   43989: out<=0;
   43990: out<=1;
   43991: out<=1;
   43992: out<=0;
   43993: out<=0;
   43994: out<=0;
   43995: out<=0;
   43996: out<=0;
   43997: out<=1;
   43998: out<=1;
   43999: out<=0;
   44000: out<=1;
   44001: out<=0;
   44002: out<=0;
   44003: out<=1;
   44004: out<=1;
   44005: out<=1;
   44006: out<=1;
   44007: out<=1;
   44008: out<=0;
   44009: out<=0;
   44010: out<=1;
   44011: out<=1;
   44012: out<=0;
   44013: out<=1;
   44014: out<=0;
   44015: out<=1;
   44016: out<=0;
   44017: out<=0;
   44018: out<=0;
   44019: out<=0;
   44020: out<=1;
   44021: out<=0;
   44022: out<=0;
   44023: out<=1;
   44024: out<=0;
   44025: out<=1;
   44026: out<=0;
   44027: out<=1;
   44028: out<=1;
   44029: out<=1;
   44030: out<=0;
   44031: out<=0;
   44032: out<=0;
   44033: out<=1;
   44034: out<=1;
   44035: out<=0;
   44036: out<=1;
   44037: out<=1;
   44038: out<=1;
   44039: out<=1;
   44040: out<=0;
   44041: out<=0;
   44042: out<=1;
   44043: out<=1;
   44044: out<=1;
   44045: out<=0;
   44046: out<=1;
   44047: out<=0;
   44048: out<=1;
   44049: out<=1;
   44050: out<=1;
   44051: out<=1;
   44052: out<=1;
   44053: out<=0;
   44054: out<=0;
   44055: out<=1;
   44056: out<=0;
   44057: out<=1;
   44058: out<=0;
   44059: out<=1;
   44060: out<=0;
   44061: out<=0;
   44062: out<=1;
   44063: out<=1;
   44064: out<=0;
   44065: out<=0;
   44066: out<=1;
   44067: out<=1;
   44068: out<=0;
   44069: out<=1;
   44070: out<=0;
   44071: out<=1;
   44072: out<=0;
   44073: out<=1;
   44074: out<=1;
   44075: out<=0;
   44076: out<=0;
   44077: out<=0;
   44078: out<=0;
   44079: out<=0;
   44080: out<=1;
   44081: out<=0;
   44082: out<=1;
   44083: out<=0;
   44084: out<=0;
   44085: out<=0;
   44086: out<=1;
   44087: out<=1;
   44088: out<=0;
   44089: out<=0;
   44090: out<=0;
   44091: out<=0;
   44092: out<=1;
   44093: out<=0;
   44094: out<=0;
   44095: out<=1;
   44096: out<=0;
   44097: out<=1;
   44098: out<=1;
   44099: out<=0;
   44100: out<=1;
   44101: out<=1;
   44102: out<=1;
   44103: out<=1;
   44104: out<=0;
   44105: out<=0;
   44106: out<=1;
   44107: out<=1;
   44108: out<=1;
   44109: out<=0;
   44110: out<=1;
   44111: out<=0;
   44112: out<=0;
   44113: out<=0;
   44114: out<=0;
   44115: out<=0;
   44116: out<=0;
   44117: out<=1;
   44118: out<=1;
   44119: out<=0;
   44120: out<=1;
   44121: out<=0;
   44122: out<=1;
   44123: out<=0;
   44124: out<=1;
   44125: out<=1;
   44126: out<=0;
   44127: out<=0;
   44128: out<=1;
   44129: out<=1;
   44130: out<=0;
   44131: out<=0;
   44132: out<=1;
   44133: out<=0;
   44134: out<=1;
   44135: out<=0;
   44136: out<=1;
   44137: out<=0;
   44138: out<=0;
   44139: out<=1;
   44140: out<=1;
   44141: out<=1;
   44142: out<=1;
   44143: out<=1;
   44144: out<=1;
   44145: out<=0;
   44146: out<=1;
   44147: out<=0;
   44148: out<=0;
   44149: out<=0;
   44150: out<=1;
   44151: out<=1;
   44152: out<=0;
   44153: out<=0;
   44154: out<=0;
   44155: out<=0;
   44156: out<=1;
   44157: out<=0;
   44158: out<=0;
   44159: out<=1;
   44160: out<=1;
   44161: out<=0;
   44162: out<=0;
   44163: out<=1;
   44164: out<=0;
   44165: out<=0;
   44166: out<=0;
   44167: out<=0;
   44168: out<=1;
   44169: out<=1;
   44170: out<=0;
   44171: out<=0;
   44172: out<=0;
   44173: out<=1;
   44174: out<=0;
   44175: out<=1;
   44176: out<=1;
   44177: out<=1;
   44178: out<=1;
   44179: out<=1;
   44180: out<=1;
   44181: out<=0;
   44182: out<=0;
   44183: out<=1;
   44184: out<=0;
   44185: out<=1;
   44186: out<=0;
   44187: out<=1;
   44188: out<=0;
   44189: out<=0;
   44190: out<=1;
   44191: out<=1;
   44192: out<=1;
   44193: out<=1;
   44194: out<=0;
   44195: out<=0;
   44196: out<=1;
   44197: out<=0;
   44198: out<=1;
   44199: out<=0;
   44200: out<=1;
   44201: out<=0;
   44202: out<=0;
   44203: out<=1;
   44204: out<=1;
   44205: out<=1;
   44206: out<=1;
   44207: out<=1;
   44208: out<=1;
   44209: out<=0;
   44210: out<=1;
   44211: out<=0;
   44212: out<=0;
   44213: out<=0;
   44214: out<=1;
   44215: out<=1;
   44216: out<=0;
   44217: out<=0;
   44218: out<=0;
   44219: out<=0;
   44220: out<=1;
   44221: out<=0;
   44222: out<=0;
   44223: out<=1;
   44224: out<=1;
   44225: out<=0;
   44226: out<=0;
   44227: out<=1;
   44228: out<=0;
   44229: out<=0;
   44230: out<=0;
   44231: out<=0;
   44232: out<=1;
   44233: out<=1;
   44234: out<=0;
   44235: out<=0;
   44236: out<=0;
   44237: out<=1;
   44238: out<=0;
   44239: out<=1;
   44240: out<=0;
   44241: out<=0;
   44242: out<=0;
   44243: out<=0;
   44244: out<=0;
   44245: out<=1;
   44246: out<=1;
   44247: out<=0;
   44248: out<=1;
   44249: out<=0;
   44250: out<=1;
   44251: out<=0;
   44252: out<=1;
   44253: out<=1;
   44254: out<=0;
   44255: out<=0;
   44256: out<=0;
   44257: out<=0;
   44258: out<=1;
   44259: out<=1;
   44260: out<=0;
   44261: out<=1;
   44262: out<=0;
   44263: out<=1;
   44264: out<=0;
   44265: out<=1;
   44266: out<=1;
   44267: out<=0;
   44268: out<=0;
   44269: out<=0;
   44270: out<=0;
   44271: out<=0;
   44272: out<=1;
   44273: out<=0;
   44274: out<=1;
   44275: out<=0;
   44276: out<=0;
   44277: out<=0;
   44278: out<=1;
   44279: out<=1;
   44280: out<=0;
   44281: out<=0;
   44282: out<=0;
   44283: out<=0;
   44284: out<=1;
   44285: out<=0;
   44286: out<=0;
   44287: out<=1;
   44288: out<=0;
   44289: out<=0;
   44290: out<=0;
   44291: out<=0;
   44292: out<=0;
   44293: out<=1;
   44294: out<=1;
   44295: out<=0;
   44296: out<=1;
   44297: out<=0;
   44298: out<=1;
   44299: out<=0;
   44300: out<=1;
   44301: out<=1;
   44302: out<=0;
   44303: out<=0;
   44304: out<=0;
   44305: out<=1;
   44306: out<=1;
   44307: out<=0;
   44308: out<=1;
   44309: out<=1;
   44310: out<=1;
   44311: out<=1;
   44312: out<=0;
   44313: out<=0;
   44314: out<=1;
   44315: out<=1;
   44316: out<=1;
   44317: out<=0;
   44318: out<=1;
   44319: out<=0;
   44320: out<=1;
   44321: out<=0;
   44322: out<=1;
   44323: out<=0;
   44324: out<=0;
   44325: out<=0;
   44326: out<=1;
   44327: out<=1;
   44328: out<=0;
   44329: out<=0;
   44330: out<=0;
   44331: out<=0;
   44332: out<=1;
   44333: out<=0;
   44334: out<=0;
   44335: out<=1;
   44336: out<=1;
   44337: out<=1;
   44338: out<=0;
   44339: out<=0;
   44340: out<=1;
   44341: out<=0;
   44342: out<=1;
   44343: out<=0;
   44344: out<=1;
   44345: out<=0;
   44346: out<=0;
   44347: out<=1;
   44348: out<=1;
   44349: out<=1;
   44350: out<=1;
   44351: out<=1;
   44352: out<=1;
   44353: out<=1;
   44354: out<=1;
   44355: out<=1;
   44356: out<=1;
   44357: out<=0;
   44358: out<=0;
   44359: out<=1;
   44360: out<=0;
   44361: out<=1;
   44362: out<=0;
   44363: out<=1;
   44364: out<=0;
   44365: out<=0;
   44366: out<=1;
   44367: out<=1;
   44368: out<=0;
   44369: out<=1;
   44370: out<=1;
   44371: out<=0;
   44372: out<=1;
   44373: out<=1;
   44374: out<=1;
   44375: out<=1;
   44376: out<=0;
   44377: out<=0;
   44378: out<=1;
   44379: out<=1;
   44380: out<=1;
   44381: out<=0;
   44382: out<=1;
   44383: out<=0;
   44384: out<=1;
   44385: out<=0;
   44386: out<=1;
   44387: out<=0;
   44388: out<=0;
   44389: out<=0;
   44390: out<=1;
   44391: out<=1;
   44392: out<=0;
   44393: out<=0;
   44394: out<=0;
   44395: out<=0;
   44396: out<=1;
   44397: out<=0;
   44398: out<=0;
   44399: out<=1;
   44400: out<=0;
   44401: out<=0;
   44402: out<=1;
   44403: out<=1;
   44404: out<=0;
   44405: out<=1;
   44406: out<=0;
   44407: out<=1;
   44408: out<=0;
   44409: out<=1;
   44410: out<=1;
   44411: out<=0;
   44412: out<=0;
   44413: out<=0;
   44414: out<=0;
   44415: out<=0;
   44416: out<=0;
   44417: out<=0;
   44418: out<=0;
   44419: out<=0;
   44420: out<=0;
   44421: out<=1;
   44422: out<=1;
   44423: out<=0;
   44424: out<=1;
   44425: out<=0;
   44426: out<=1;
   44427: out<=0;
   44428: out<=1;
   44429: out<=1;
   44430: out<=0;
   44431: out<=0;
   44432: out<=1;
   44433: out<=0;
   44434: out<=0;
   44435: out<=1;
   44436: out<=0;
   44437: out<=0;
   44438: out<=0;
   44439: out<=0;
   44440: out<=1;
   44441: out<=1;
   44442: out<=0;
   44443: out<=0;
   44444: out<=0;
   44445: out<=1;
   44446: out<=0;
   44447: out<=1;
   44448: out<=1;
   44449: out<=0;
   44450: out<=1;
   44451: out<=0;
   44452: out<=0;
   44453: out<=0;
   44454: out<=1;
   44455: out<=1;
   44456: out<=0;
   44457: out<=0;
   44458: out<=0;
   44459: out<=0;
   44460: out<=1;
   44461: out<=0;
   44462: out<=0;
   44463: out<=1;
   44464: out<=0;
   44465: out<=0;
   44466: out<=1;
   44467: out<=1;
   44468: out<=0;
   44469: out<=1;
   44470: out<=0;
   44471: out<=1;
   44472: out<=0;
   44473: out<=1;
   44474: out<=1;
   44475: out<=0;
   44476: out<=0;
   44477: out<=0;
   44478: out<=0;
   44479: out<=0;
   44480: out<=1;
   44481: out<=1;
   44482: out<=1;
   44483: out<=1;
   44484: out<=1;
   44485: out<=0;
   44486: out<=0;
   44487: out<=1;
   44488: out<=0;
   44489: out<=1;
   44490: out<=0;
   44491: out<=1;
   44492: out<=0;
   44493: out<=0;
   44494: out<=1;
   44495: out<=1;
   44496: out<=1;
   44497: out<=0;
   44498: out<=0;
   44499: out<=1;
   44500: out<=0;
   44501: out<=0;
   44502: out<=0;
   44503: out<=0;
   44504: out<=1;
   44505: out<=1;
   44506: out<=0;
   44507: out<=0;
   44508: out<=0;
   44509: out<=1;
   44510: out<=0;
   44511: out<=1;
   44512: out<=1;
   44513: out<=0;
   44514: out<=1;
   44515: out<=0;
   44516: out<=0;
   44517: out<=0;
   44518: out<=1;
   44519: out<=1;
   44520: out<=0;
   44521: out<=0;
   44522: out<=0;
   44523: out<=0;
   44524: out<=1;
   44525: out<=0;
   44526: out<=0;
   44527: out<=1;
   44528: out<=1;
   44529: out<=1;
   44530: out<=0;
   44531: out<=0;
   44532: out<=1;
   44533: out<=0;
   44534: out<=1;
   44535: out<=0;
   44536: out<=1;
   44537: out<=0;
   44538: out<=0;
   44539: out<=1;
   44540: out<=1;
   44541: out<=1;
   44542: out<=1;
   44543: out<=1;
   44544: out<=1;
   44545: out<=1;
   44546: out<=0;
   44547: out<=0;
   44548: out<=1;
   44549: out<=0;
   44550: out<=1;
   44551: out<=0;
   44552: out<=1;
   44553: out<=0;
   44554: out<=0;
   44555: out<=1;
   44556: out<=1;
   44557: out<=1;
   44558: out<=1;
   44559: out<=1;
   44560: out<=1;
   44561: out<=0;
   44562: out<=1;
   44563: out<=0;
   44564: out<=0;
   44565: out<=0;
   44566: out<=1;
   44567: out<=1;
   44568: out<=0;
   44569: out<=0;
   44570: out<=0;
   44571: out<=0;
   44572: out<=1;
   44573: out<=0;
   44574: out<=0;
   44575: out<=1;
   44576: out<=1;
   44577: out<=0;
   44578: out<=0;
   44579: out<=1;
   44580: out<=0;
   44581: out<=0;
   44582: out<=0;
   44583: out<=0;
   44584: out<=1;
   44585: out<=1;
   44586: out<=0;
   44587: out<=0;
   44588: out<=0;
   44589: out<=1;
   44590: out<=0;
   44591: out<=1;
   44592: out<=1;
   44593: out<=1;
   44594: out<=1;
   44595: out<=1;
   44596: out<=1;
   44597: out<=0;
   44598: out<=0;
   44599: out<=1;
   44600: out<=0;
   44601: out<=1;
   44602: out<=0;
   44603: out<=1;
   44604: out<=0;
   44605: out<=0;
   44606: out<=1;
   44607: out<=1;
   44608: out<=0;
   44609: out<=0;
   44610: out<=1;
   44611: out<=1;
   44612: out<=0;
   44613: out<=1;
   44614: out<=0;
   44615: out<=1;
   44616: out<=0;
   44617: out<=1;
   44618: out<=1;
   44619: out<=0;
   44620: out<=0;
   44621: out<=0;
   44622: out<=0;
   44623: out<=0;
   44624: out<=1;
   44625: out<=0;
   44626: out<=1;
   44627: out<=0;
   44628: out<=0;
   44629: out<=0;
   44630: out<=1;
   44631: out<=1;
   44632: out<=0;
   44633: out<=0;
   44634: out<=0;
   44635: out<=0;
   44636: out<=1;
   44637: out<=0;
   44638: out<=0;
   44639: out<=1;
   44640: out<=1;
   44641: out<=0;
   44642: out<=0;
   44643: out<=1;
   44644: out<=0;
   44645: out<=0;
   44646: out<=0;
   44647: out<=0;
   44648: out<=1;
   44649: out<=1;
   44650: out<=0;
   44651: out<=0;
   44652: out<=0;
   44653: out<=1;
   44654: out<=0;
   44655: out<=1;
   44656: out<=0;
   44657: out<=0;
   44658: out<=0;
   44659: out<=0;
   44660: out<=0;
   44661: out<=1;
   44662: out<=1;
   44663: out<=0;
   44664: out<=1;
   44665: out<=0;
   44666: out<=1;
   44667: out<=0;
   44668: out<=1;
   44669: out<=1;
   44670: out<=0;
   44671: out<=0;
   44672: out<=0;
   44673: out<=0;
   44674: out<=1;
   44675: out<=1;
   44676: out<=0;
   44677: out<=1;
   44678: out<=0;
   44679: out<=1;
   44680: out<=0;
   44681: out<=1;
   44682: out<=1;
   44683: out<=0;
   44684: out<=0;
   44685: out<=0;
   44686: out<=0;
   44687: out<=0;
   44688: out<=1;
   44689: out<=0;
   44690: out<=1;
   44691: out<=0;
   44692: out<=0;
   44693: out<=0;
   44694: out<=1;
   44695: out<=1;
   44696: out<=0;
   44697: out<=0;
   44698: out<=0;
   44699: out<=0;
   44700: out<=1;
   44701: out<=0;
   44702: out<=0;
   44703: out<=1;
   44704: out<=0;
   44705: out<=1;
   44706: out<=1;
   44707: out<=0;
   44708: out<=1;
   44709: out<=1;
   44710: out<=1;
   44711: out<=1;
   44712: out<=0;
   44713: out<=0;
   44714: out<=1;
   44715: out<=1;
   44716: out<=1;
   44717: out<=0;
   44718: out<=1;
   44719: out<=0;
   44720: out<=1;
   44721: out<=1;
   44722: out<=1;
   44723: out<=1;
   44724: out<=1;
   44725: out<=0;
   44726: out<=0;
   44727: out<=1;
   44728: out<=0;
   44729: out<=1;
   44730: out<=0;
   44731: out<=1;
   44732: out<=0;
   44733: out<=0;
   44734: out<=1;
   44735: out<=1;
   44736: out<=1;
   44737: out<=1;
   44738: out<=0;
   44739: out<=0;
   44740: out<=1;
   44741: out<=0;
   44742: out<=1;
   44743: out<=0;
   44744: out<=1;
   44745: out<=0;
   44746: out<=0;
   44747: out<=1;
   44748: out<=1;
   44749: out<=1;
   44750: out<=1;
   44751: out<=1;
   44752: out<=1;
   44753: out<=0;
   44754: out<=1;
   44755: out<=0;
   44756: out<=0;
   44757: out<=0;
   44758: out<=1;
   44759: out<=1;
   44760: out<=0;
   44761: out<=0;
   44762: out<=0;
   44763: out<=0;
   44764: out<=1;
   44765: out<=0;
   44766: out<=0;
   44767: out<=1;
   44768: out<=0;
   44769: out<=1;
   44770: out<=1;
   44771: out<=0;
   44772: out<=1;
   44773: out<=1;
   44774: out<=1;
   44775: out<=1;
   44776: out<=0;
   44777: out<=0;
   44778: out<=1;
   44779: out<=1;
   44780: out<=1;
   44781: out<=0;
   44782: out<=1;
   44783: out<=0;
   44784: out<=0;
   44785: out<=0;
   44786: out<=0;
   44787: out<=0;
   44788: out<=0;
   44789: out<=1;
   44790: out<=1;
   44791: out<=0;
   44792: out<=1;
   44793: out<=0;
   44794: out<=1;
   44795: out<=0;
   44796: out<=1;
   44797: out<=1;
   44798: out<=0;
   44799: out<=0;
   44800: out<=1;
   44801: out<=0;
   44802: out<=1;
   44803: out<=0;
   44804: out<=0;
   44805: out<=0;
   44806: out<=1;
   44807: out<=1;
   44808: out<=0;
   44809: out<=0;
   44810: out<=0;
   44811: out<=0;
   44812: out<=1;
   44813: out<=0;
   44814: out<=0;
   44815: out<=1;
   44816: out<=0;
   44817: out<=0;
   44818: out<=1;
   44819: out<=1;
   44820: out<=0;
   44821: out<=1;
   44822: out<=0;
   44823: out<=1;
   44824: out<=0;
   44825: out<=1;
   44826: out<=1;
   44827: out<=0;
   44828: out<=0;
   44829: out<=0;
   44830: out<=0;
   44831: out<=0;
   44832: out<=0;
   44833: out<=0;
   44834: out<=0;
   44835: out<=0;
   44836: out<=0;
   44837: out<=1;
   44838: out<=1;
   44839: out<=0;
   44840: out<=1;
   44841: out<=0;
   44842: out<=1;
   44843: out<=0;
   44844: out<=1;
   44845: out<=1;
   44846: out<=0;
   44847: out<=0;
   44848: out<=1;
   44849: out<=0;
   44850: out<=0;
   44851: out<=1;
   44852: out<=0;
   44853: out<=0;
   44854: out<=0;
   44855: out<=0;
   44856: out<=1;
   44857: out<=1;
   44858: out<=0;
   44859: out<=0;
   44860: out<=0;
   44861: out<=1;
   44862: out<=0;
   44863: out<=1;
   44864: out<=1;
   44865: out<=0;
   44866: out<=1;
   44867: out<=0;
   44868: out<=0;
   44869: out<=0;
   44870: out<=1;
   44871: out<=1;
   44872: out<=0;
   44873: out<=0;
   44874: out<=0;
   44875: out<=0;
   44876: out<=1;
   44877: out<=0;
   44878: out<=0;
   44879: out<=1;
   44880: out<=1;
   44881: out<=1;
   44882: out<=0;
   44883: out<=0;
   44884: out<=1;
   44885: out<=0;
   44886: out<=1;
   44887: out<=0;
   44888: out<=1;
   44889: out<=0;
   44890: out<=0;
   44891: out<=1;
   44892: out<=1;
   44893: out<=1;
   44894: out<=1;
   44895: out<=1;
   44896: out<=1;
   44897: out<=1;
   44898: out<=1;
   44899: out<=1;
   44900: out<=1;
   44901: out<=0;
   44902: out<=0;
   44903: out<=1;
   44904: out<=0;
   44905: out<=1;
   44906: out<=0;
   44907: out<=1;
   44908: out<=0;
   44909: out<=0;
   44910: out<=1;
   44911: out<=1;
   44912: out<=1;
   44913: out<=0;
   44914: out<=0;
   44915: out<=1;
   44916: out<=0;
   44917: out<=0;
   44918: out<=0;
   44919: out<=0;
   44920: out<=1;
   44921: out<=1;
   44922: out<=0;
   44923: out<=0;
   44924: out<=0;
   44925: out<=1;
   44926: out<=0;
   44927: out<=1;
   44928: out<=1;
   44929: out<=0;
   44930: out<=1;
   44931: out<=0;
   44932: out<=0;
   44933: out<=0;
   44934: out<=1;
   44935: out<=1;
   44936: out<=0;
   44937: out<=0;
   44938: out<=0;
   44939: out<=0;
   44940: out<=1;
   44941: out<=0;
   44942: out<=0;
   44943: out<=1;
   44944: out<=1;
   44945: out<=1;
   44946: out<=0;
   44947: out<=0;
   44948: out<=1;
   44949: out<=0;
   44950: out<=1;
   44951: out<=0;
   44952: out<=1;
   44953: out<=0;
   44954: out<=0;
   44955: out<=1;
   44956: out<=1;
   44957: out<=1;
   44958: out<=1;
   44959: out<=1;
   44960: out<=0;
   44961: out<=0;
   44962: out<=0;
   44963: out<=0;
   44964: out<=0;
   44965: out<=1;
   44966: out<=1;
   44967: out<=0;
   44968: out<=1;
   44969: out<=0;
   44970: out<=1;
   44971: out<=0;
   44972: out<=1;
   44973: out<=1;
   44974: out<=0;
   44975: out<=0;
   44976: out<=0;
   44977: out<=1;
   44978: out<=1;
   44979: out<=0;
   44980: out<=1;
   44981: out<=1;
   44982: out<=1;
   44983: out<=1;
   44984: out<=0;
   44985: out<=0;
   44986: out<=1;
   44987: out<=1;
   44988: out<=1;
   44989: out<=0;
   44990: out<=1;
   44991: out<=0;
   44992: out<=1;
   44993: out<=0;
   44994: out<=1;
   44995: out<=0;
   44996: out<=0;
   44997: out<=0;
   44998: out<=1;
   44999: out<=1;
   45000: out<=0;
   45001: out<=0;
   45002: out<=0;
   45003: out<=0;
   45004: out<=1;
   45005: out<=0;
   45006: out<=0;
   45007: out<=1;
   45008: out<=0;
   45009: out<=0;
   45010: out<=1;
   45011: out<=1;
   45012: out<=0;
   45013: out<=1;
   45014: out<=0;
   45015: out<=1;
   45016: out<=0;
   45017: out<=1;
   45018: out<=1;
   45019: out<=0;
   45020: out<=0;
   45021: out<=0;
   45022: out<=0;
   45023: out<=0;
   45024: out<=1;
   45025: out<=1;
   45026: out<=1;
   45027: out<=1;
   45028: out<=1;
   45029: out<=0;
   45030: out<=0;
   45031: out<=1;
   45032: out<=0;
   45033: out<=1;
   45034: out<=0;
   45035: out<=1;
   45036: out<=0;
   45037: out<=0;
   45038: out<=1;
   45039: out<=1;
   45040: out<=0;
   45041: out<=1;
   45042: out<=1;
   45043: out<=0;
   45044: out<=1;
   45045: out<=1;
   45046: out<=1;
   45047: out<=1;
   45048: out<=0;
   45049: out<=0;
   45050: out<=1;
   45051: out<=1;
   45052: out<=1;
   45053: out<=0;
   45054: out<=1;
   45055: out<=0;
   45056: out<=0;
   45057: out<=1;
   45058: out<=0;
   45059: out<=1;
   45060: out<=0;
   45061: out<=0;
   45062: out<=1;
   45063: out<=1;
   45064: out<=1;
   45065: out<=1;
   45066: out<=1;
   45067: out<=1;
   45068: out<=1;
   45069: out<=0;
   45070: out<=0;
   45071: out<=1;
   45072: out<=1;
   45073: out<=1;
   45074: out<=0;
   45075: out<=0;
   45076: out<=0;
   45077: out<=1;
   45078: out<=0;
   45079: out<=1;
   45080: out<=1;
   45081: out<=0;
   45082: out<=0;
   45083: out<=1;
   45084: out<=0;
   45085: out<=0;
   45086: out<=0;
   45087: out<=0;
   45088: out<=0;
   45089: out<=0;
   45090: out<=0;
   45091: out<=0;
   45092: out<=1;
   45093: out<=0;
   45094: out<=0;
   45095: out<=1;
   45096: out<=1;
   45097: out<=0;
   45098: out<=1;
   45099: out<=0;
   45100: out<=0;
   45101: out<=0;
   45102: out<=1;
   45103: out<=1;
   45104: out<=1;
   45105: out<=0;
   45106: out<=0;
   45107: out<=1;
   45108: out<=1;
   45109: out<=1;
   45110: out<=1;
   45111: out<=1;
   45112: out<=1;
   45113: out<=1;
   45114: out<=0;
   45115: out<=0;
   45116: out<=1;
   45117: out<=0;
   45118: out<=1;
   45119: out<=0;
   45120: out<=0;
   45121: out<=1;
   45122: out<=0;
   45123: out<=1;
   45124: out<=0;
   45125: out<=0;
   45126: out<=1;
   45127: out<=1;
   45128: out<=1;
   45129: out<=1;
   45130: out<=1;
   45131: out<=1;
   45132: out<=1;
   45133: out<=0;
   45134: out<=0;
   45135: out<=1;
   45136: out<=0;
   45137: out<=0;
   45138: out<=1;
   45139: out<=1;
   45140: out<=1;
   45141: out<=0;
   45142: out<=1;
   45143: out<=0;
   45144: out<=0;
   45145: out<=1;
   45146: out<=1;
   45147: out<=0;
   45148: out<=1;
   45149: out<=1;
   45150: out<=1;
   45151: out<=1;
   45152: out<=1;
   45153: out<=1;
   45154: out<=1;
   45155: out<=1;
   45156: out<=0;
   45157: out<=1;
   45158: out<=1;
   45159: out<=0;
   45160: out<=0;
   45161: out<=1;
   45162: out<=0;
   45163: out<=1;
   45164: out<=1;
   45165: out<=1;
   45166: out<=0;
   45167: out<=0;
   45168: out<=1;
   45169: out<=0;
   45170: out<=0;
   45171: out<=1;
   45172: out<=1;
   45173: out<=1;
   45174: out<=1;
   45175: out<=1;
   45176: out<=1;
   45177: out<=1;
   45178: out<=0;
   45179: out<=0;
   45180: out<=1;
   45181: out<=0;
   45182: out<=1;
   45183: out<=0;
   45184: out<=0;
   45185: out<=1;
   45186: out<=0;
   45187: out<=1;
   45188: out<=0;
   45189: out<=0;
   45190: out<=1;
   45191: out<=1;
   45192: out<=1;
   45193: out<=1;
   45194: out<=1;
   45195: out<=1;
   45196: out<=1;
   45197: out<=0;
   45198: out<=0;
   45199: out<=1;
   45200: out<=0;
   45201: out<=0;
   45202: out<=1;
   45203: out<=1;
   45204: out<=1;
   45205: out<=0;
   45206: out<=1;
   45207: out<=0;
   45208: out<=0;
   45209: out<=1;
   45210: out<=1;
   45211: out<=0;
   45212: out<=1;
   45213: out<=1;
   45214: out<=1;
   45215: out<=1;
   45216: out<=0;
   45217: out<=0;
   45218: out<=0;
   45219: out<=0;
   45220: out<=1;
   45221: out<=0;
   45222: out<=0;
   45223: out<=1;
   45224: out<=1;
   45225: out<=0;
   45226: out<=1;
   45227: out<=0;
   45228: out<=0;
   45229: out<=0;
   45230: out<=1;
   45231: out<=1;
   45232: out<=0;
   45233: out<=1;
   45234: out<=1;
   45235: out<=0;
   45236: out<=0;
   45237: out<=0;
   45238: out<=0;
   45239: out<=0;
   45240: out<=0;
   45241: out<=0;
   45242: out<=1;
   45243: out<=1;
   45244: out<=0;
   45245: out<=1;
   45246: out<=0;
   45247: out<=1;
   45248: out<=0;
   45249: out<=1;
   45250: out<=0;
   45251: out<=1;
   45252: out<=0;
   45253: out<=0;
   45254: out<=1;
   45255: out<=1;
   45256: out<=1;
   45257: out<=1;
   45258: out<=1;
   45259: out<=1;
   45260: out<=1;
   45261: out<=0;
   45262: out<=0;
   45263: out<=1;
   45264: out<=1;
   45265: out<=1;
   45266: out<=0;
   45267: out<=0;
   45268: out<=0;
   45269: out<=1;
   45270: out<=0;
   45271: out<=1;
   45272: out<=1;
   45273: out<=0;
   45274: out<=0;
   45275: out<=1;
   45276: out<=0;
   45277: out<=0;
   45278: out<=0;
   45279: out<=0;
   45280: out<=1;
   45281: out<=1;
   45282: out<=1;
   45283: out<=1;
   45284: out<=0;
   45285: out<=1;
   45286: out<=1;
   45287: out<=0;
   45288: out<=0;
   45289: out<=1;
   45290: out<=0;
   45291: out<=1;
   45292: out<=1;
   45293: out<=1;
   45294: out<=0;
   45295: out<=0;
   45296: out<=0;
   45297: out<=1;
   45298: out<=1;
   45299: out<=0;
   45300: out<=0;
   45301: out<=0;
   45302: out<=0;
   45303: out<=0;
   45304: out<=0;
   45305: out<=0;
   45306: out<=1;
   45307: out<=1;
   45308: out<=0;
   45309: out<=1;
   45310: out<=0;
   45311: out<=1;
   45312: out<=0;
   45313: out<=0;
   45314: out<=1;
   45315: out<=1;
   45316: out<=1;
   45317: out<=0;
   45318: out<=1;
   45319: out<=0;
   45320: out<=0;
   45321: out<=1;
   45322: out<=1;
   45323: out<=0;
   45324: out<=1;
   45325: out<=1;
   45326: out<=1;
   45327: out<=1;
   45328: out<=0;
   45329: out<=1;
   45330: out<=0;
   45331: out<=1;
   45332: out<=0;
   45333: out<=0;
   45334: out<=1;
   45335: out<=1;
   45336: out<=1;
   45337: out<=1;
   45338: out<=1;
   45339: out<=1;
   45340: out<=1;
   45341: out<=0;
   45342: out<=0;
   45343: out<=1;
   45344: out<=1;
   45345: out<=0;
   45346: out<=0;
   45347: out<=1;
   45348: out<=1;
   45349: out<=1;
   45350: out<=1;
   45351: out<=1;
   45352: out<=1;
   45353: out<=1;
   45354: out<=0;
   45355: out<=0;
   45356: out<=1;
   45357: out<=0;
   45358: out<=1;
   45359: out<=0;
   45360: out<=1;
   45361: out<=1;
   45362: out<=1;
   45363: out<=1;
   45364: out<=0;
   45365: out<=1;
   45366: out<=1;
   45367: out<=0;
   45368: out<=0;
   45369: out<=1;
   45370: out<=0;
   45371: out<=1;
   45372: out<=1;
   45373: out<=1;
   45374: out<=0;
   45375: out<=0;
   45376: out<=1;
   45377: out<=1;
   45378: out<=0;
   45379: out<=0;
   45380: out<=0;
   45381: out<=1;
   45382: out<=0;
   45383: out<=1;
   45384: out<=1;
   45385: out<=0;
   45386: out<=0;
   45387: out<=1;
   45388: out<=0;
   45389: out<=0;
   45390: out<=0;
   45391: out<=0;
   45392: out<=0;
   45393: out<=1;
   45394: out<=0;
   45395: out<=1;
   45396: out<=0;
   45397: out<=0;
   45398: out<=1;
   45399: out<=1;
   45400: out<=1;
   45401: out<=1;
   45402: out<=1;
   45403: out<=1;
   45404: out<=1;
   45405: out<=0;
   45406: out<=0;
   45407: out<=1;
   45408: out<=1;
   45409: out<=0;
   45410: out<=0;
   45411: out<=1;
   45412: out<=1;
   45413: out<=1;
   45414: out<=1;
   45415: out<=1;
   45416: out<=1;
   45417: out<=1;
   45418: out<=0;
   45419: out<=0;
   45420: out<=1;
   45421: out<=0;
   45422: out<=1;
   45423: out<=0;
   45424: out<=0;
   45425: out<=0;
   45426: out<=0;
   45427: out<=0;
   45428: out<=1;
   45429: out<=0;
   45430: out<=0;
   45431: out<=1;
   45432: out<=1;
   45433: out<=0;
   45434: out<=1;
   45435: out<=0;
   45436: out<=0;
   45437: out<=0;
   45438: out<=1;
   45439: out<=1;
   45440: out<=1;
   45441: out<=1;
   45442: out<=0;
   45443: out<=0;
   45444: out<=0;
   45445: out<=1;
   45446: out<=0;
   45447: out<=1;
   45448: out<=1;
   45449: out<=0;
   45450: out<=0;
   45451: out<=1;
   45452: out<=0;
   45453: out<=0;
   45454: out<=0;
   45455: out<=0;
   45456: out<=0;
   45457: out<=1;
   45458: out<=0;
   45459: out<=1;
   45460: out<=0;
   45461: out<=0;
   45462: out<=1;
   45463: out<=1;
   45464: out<=1;
   45465: out<=1;
   45466: out<=1;
   45467: out<=1;
   45468: out<=1;
   45469: out<=0;
   45470: out<=0;
   45471: out<=1;
   45472: out<=0;
   45473: out<=1;
   45474: out<=1;
   45475: out<=0;
   45476: out<=0;
   45477: out<=0;
   45478: out<=0;
   45479: out<=0;
   45480: out<=0;
   45481: out<=0;
   45482: out<=1;
   45483: out<=1;
   45484: out<=0;
   45485: out<=1;
   45486: out<=0;
   45487: out<=1;
   45488: out<=1;
   45489: out<=1;
   45490: out<=1;
   45491: out<=1;
   45492: out<=0;
   45493: out<=1;
   45494: out<=1;
   45495: out<=0;
   45496: out<=0;
   45497: out<=1;
   45498: out<=0;
   45499: out<=1;
   45500: out<=1;
   45501: out<=1;
   45502: out<=0;
   45503: out<=0;
   45504: out<=0;
   45505: out<=0;
   45506: out<=1;
   45507: out<=1;
   45508: out<=1;
   45509: out<=0;
   45510: out<=1;
   45511: out<=0;
   45512: out<=0;
   45513: out<=1;
   45514: out<=1;
   45515: out<=0;
   45516: out<=1;
   45517: out<=1;
   45518: out<=1;
   45519: out<=1;
   45520: out<=0;
   45521: out<=1;
   45522: out<=0;
   45523: out<=1;
   45524: out<=0;
   45525: out<=0;
   45526: out<=1;
   45527: out<=1;
   45528: out<=1;
   45529: out<=1;
   45530: out<=1;
   45531: out<=1;
   45532: out<=1;
   45533: out<=0;
   45534: out<=0;
   45535: out<=1;
   45536: out<=0;
   45537: out<=1;
   45538: out<=1;
   45539: out<=0;
   45540: out<=0;
   45541: out<=0;
   45542: out<=0;
   45543: out<=0;
   45544: out<=0;
   45545: out<=0;
   45546: out<=1;
   45547: out<=1;
   45548: out<=0;
   45549: out<=1;
   45550: out<=0;
   45551: out<=1;
   45552: out<=0;
   45553: out<=0;
   45554: out<=0;
   45555: out<=0;
   45556: out<=1;
   45557: out<=0;
   45558: out<=0;
   45559: out<=1;
   45560: out<=1;
   45561: out<=0;
   45562: out<=1;
   45563: out<=0;
   45564: out<=0;
   45565: out<=0;
   45566: out<=1;
   45567: out<=1;
   45568: out<=0;
   45569: out<=0;
   45570: out<=0;
   45571: out<=0;
   45572: out<=1;
   45573: out<=0;
   45574: out<=0;
   45575: out<=1;
   45576: out<=1;
   45577: out<=0;
   45578: out<=1;
   45579: out<=0;
   45580: out<=0;
   45581: out<=0;
   45582: out<=1;
   45583: out<=1;
   45584: out<=0;
   45585: out<=1;
   45586: out<=1;
   45587: out<=0;
   45588: out<=0;
   45589: out<=0;
   45590: out<=0;
   45591: out<=0;
   45592: out<=0;
   45593: out<=0;
   45594: out<=1;
   45595: out<=1;
   45596: out<=0;
   45597: out<=1;
   45598: out<=0;
   45599: out<=1;
   45600: out<=0;
   45601: out<=1;
   45602: out<=0;
   45603: out<=1;
   45604: out<=0;
   45605: out<=0;
   45606: out<=1;
   45607: out<=1;
   45608: out<=1;
   45609: out<=1;
   45610: out<=1;
   45611: out<=1;
   45612: out<=1;
   45613: out<=0;
   45614: out<=0;
   45615: out<=1;
   45616: out<=0;
   45617: out<=0;
   45618: out<=1;
   45619: out<=1;
   45620: out<=1;
   45621: out<=0;
   45622: out<=1;
   45623: out<=0;
   45624: out<=0;
   45625: out<=1;
   45626: out<=1;
   45627: out<=0;
   45628: out<=1;
   45629: out<=1;
   45630: out<=1;
   45631: out<=1;
   45632: out<=1;
   45633: out<=1;
   45634: out<=1;
   45635: out<=1;
   45636: out<=0;
   45637: out<=1;
   45638: out<=1;
   45639: out<=0;
   45640: out<=0;
   45641: out<=1;
   45642: out<=0;
   45643: out<=1;
   45644: out<=1;
   45645: out<=1;
   45646: out<=0;
   45647: out<=0;
   45648: out<=0;
   45649: out<=1;
   45650: out<=1;
   45651: out<=0;
   45652: out<=0;
   45653: out<=0;
   45654: out<=0;
   45655: out<=0;
   45656: out<=0;
   45657: out<=0;
   45658: out<=1;
   45659: out<=1;
   45660: out<=0;
   45661: out<=1;
   45662: out<=0;
   45663: out<=1;
   45664: out<=0;
   45665: out<=1;
   45666: out<=0;
   45667: out<=1;
   45668: out<=0;
   45669: out<=0;
   45670: out<=1;
   45671: out<=1;
   45672: out<=1;
   45673: out<=1;
   45674: out<=1;
   45675: out<=1;
   45676: out<=1;
   45677: out<=0;
   45678: out<=0;
   45679: out<=1;
   45680: out<=1;
   45681: out<=1;
   45682: out<=0;
   45683: out<=0;
   45684: out<=0;
   45685: out<=1;
   45686: out<=0;
   45687: out<=1;
   45688: out<=1;
   45689: out<=0;
   45690: out<=0;
   45691: out<=1;
   45692: out<=0;
   45693: out<=0;
   45694: out<=0;
   45695: out<=0;
   45696: out<=0;
   45697: out<=0;
   45698: out<=0;
   45699: out<=0;
   45700: out<=1;
   45701: out<=0;
   45702: out<=0;
   45703: out<=1;
   45704: out<=1;
   45705: out<=0;
   45706: out<=1;
   45707: out<=0;
   45708: out<=0;
   45709: out<=0;
   45710: out<=1;
   45711: out<=1;
   45712: out<=1;
   45713: out<=0;
   45714: out<=0;
   45715: out<=1;
   45716: out<=1;
   45717: out<=1;
   45718: out<=1;
   45719: out<=1;
   45720: out<=1;
   45721: out<=1;
   45722: out<=0;
   45723: out<=0;
   45724: out<=1;
   45725: out<=0;
   45726: out<=1;
   45727: out<=0;
   45728: out<=0;
   45729: out<=1;
   45730: out<=0;
   45731: out<=1;
   45732: out<=0;
   45733: out<=0;
   45734: out<=1;
   45735: out<=1;
   45736: out<=1;
   45737: out<=1;
   45738: out<=1;
   45739: out<=1;
   45740: out<=1;
   45741: out<=0;
   45742: out<=0;
   45743: out<=1;
   45744: out<=1;
   45745: out<=1;
   45746: out<=0;
   45747: out<=0;
   45748: out<=0;
   45749: out<=1;
   45750: out<=0;
   45751: out<=1;
   45752: out<=1;
   45753: out<=0;
   45754: out<=0;
   45755: out<=1;
   45756: out<=0;
   45757: out<=0;
   45758: out<=0;
   45759: out<=0;
   45760: out<=1;
   45761: out<=1;
   45762: out<=1;
   45763: out<=1;
   45764: out<=0;
   45765: out<=1;
   45766: out<=1;
   45767: out<=0;
   45768: out<=0;
   45769: out<=1;
   45770: out<=0;
   45771: out<=1;
   45772: out<=1;
   45773: out<=1;
   45774: out<=0;
   45775: out<=0;
   45776: out<=1;
   45777: out<=0;
   45778: out<=0;
   45779: out<=1;
   45780: out<=1;
   45781: out<=1;
   45782: out<=1;
   45783: out<=1;
   45784: out<=1;
   45785: out<=1;
   45786: out<=0;
   45787: out<=0;
   45788: out<=1;
   45789: out<=0;
   45790: out<=1;
   45791: out<=0;
   45792: out<=0;
   45793: out<=1;
   45794: out<=0;
   45795: out<=1;
   45796: out<=0;
   45797: out<=0;
   45798: out<=1;
   45799: out<=1;
   45800: out<=1;
   45801: out<=1;
   45802: out<=1;
   45803: out<=1;
   45804: out<=1;
   45805: out<=0;
   45806: out<=0;
   45807: out<=1;
   45808: out<=0;
   45809: out<=0;
   45810: out<=1;
   45811: out<=1;
   45812: out<=1;
   45813: out<=0;
   45814: out<=1;
   45815: out<=0;
   45816: out<=0;
   45817: out<=1;
   45818: out<=1;
   45819: out<=0;
   45820: out<=1;
   45821: out<=1;
   45822: out<=1;
   45823: out<=1;
   45824: out<=0;
   45825: out<=1;
   45826: out<=1;
   45827: out<=0;
   45828: out<=0;
   45829: out<=0;
   45830: out<=0;
   45831: out<=0;
   45832: out<=0;
   45833: out<=0;
   45834: out<=1;
   45835: out<=1;
   45836: out<=0;
   45837: out<=1;
   45838: out<=0;
   45839: out<=1;
   45840: out<=1;
   45841: out<=1;
   45842: out<=1;
   45843: out<=1;
   45844: out<=0;
   45845: out<=1;
   45846: out<=1;
   45847: out<=0;
   45848: out<=0;
   45849: out<=1;
   45850: out<=0;
   45851: out<=1;
   45852: out<=1;
   45853: out<=1;
   45854: out<=0;
   45855: out<=0;
   45856: out<=1;
   45857: out<=1;
   45858: out<=0;
   45859: out<=0;
   45860: out<=0;
   45861: out<=1;
   45862: out<=0;
   45863: out<=1;
   45864: out<=1;
   45865: out<=0;
   45866: out<=0;
   45867: out<=1;
   45868: out<=0;
   45869: out<=0;
   45870: out<=0;
   45871: out<=0;
   45872: out<=0;
   45873: out<=1;
   45874: out<=0;
   45875: out<=1;
   45876: out<=0;
   45877: out<=0;
   45878: out<=1;
   45879: out<=1;
   45880: out<=1;
   45881: out<=1;
   45882: out<=1;
   45883: out<=1;
   45884: out<=1;
   45885: out<=0;
   45886: out<=0;
   45887: out<=1;
   45888: out<=0;
   45889: out<=1;
   45890: out<=1;
   45891: out<=0;
   45892: out<=0;
   45893: out<=0;
   45894: out<=0;
   45895: out<=0;
   45896: out<=0;
   45897: out<=0;
   45898: out<=1;
   45899: out<=1;
   45900: out<=0;
   45901: out<=1;
   45902: out<=0;
   45903: out<=1;
   45904: out<=0;
   45905: out<=0;
   45906: out<=0;
   45907: out<=0;
   45908: out<=1;
   45909: out<=0;
   45910: out<=0;
   45911: out<=1;
   45912: out<=1;
   45913: out<=0;
   45914: out<=1;
   45915: out<=0;
   45916: out<=0;
   45917: out<=0;
   45918: out<=1;
   45919: out<=1;
   45920: out<=0;
   45921: out<=0;
   45922: out<=1;
   45923: out<=1;
   45924: out<=1;
   45925: out<=0;
   45926: out<=1;
   45927: out<=0;
   45928: out<=0;
   45929: out<=1;
   45930: out<=1;
   45931: out<=0;
   45932: out<=1;
   45933: out<=1;
   45934: out<=1;
   45935: out<=1;
   45936: out<=0;
   45937: out<=1;
   45938: out<=0;
   45939: out<=1;
   45940: out<=0;
   45941: out<=0;
   45942: out<=1;
   45943: out<=1;
   45944: out<=1;
   45945: out<=1;
   45946: out<=1;
   45947: out<=1;
   45948: out<=1;
   45949: out<=0;
   45950: out<=0;
   45951: out<=1;
   45952: out<=1;
   45953: out<=0;
   45954: out<=0;
   45955: out<=1;
   45956: out<=1;
   45957: out<=1;
   45958: out<=1;
   45959: out<=1;
   45960: out<=1;
   45961: out<=1;
   45962: out<=0;
   45963: out<=0;
   45964: out<=1;
   45965: out<=0;
   45966: out<=1;
   45967: out<=0;
   45968: out<=1;
   45969: out<=1;
   45970: out<=1;
   45971: out<=1;
   45972: out<=0;
   45973: out<=1;
   45974: out<=1;
   45975: out<=0;
   45976: out<=0;
   45977: out<=1;
   45978: out<=0;
   45979: out<=1;
   45980: out<=1;
   45981: out<=1;
   45982: out<=0;
   45983: out<=0;
   45984: out<=0;
   45985: out<=0;
   45986: out<=1;
   45987: out<=1;
   45988: out<=1;
   45989: out<=0;
   45990: out<=1;
   45991: out<=0;
   45992: out<=0;
   45993: out<=1;
   45994: out<=1;
   45995: out<=0;
   45996: out<=1;
   45997: out<=1;
   45998: out<=1;
   45999: out<=1;
   46000: out<=0;
   46001: out<=1;
   46002: out<=0;
   46003: out<=1;
   46004: out<=0;
   46005: out<=0;
   46006: out<=1;
   46007: out<=1;
   46008: out<=1;
   46009: out<=1;
   46010: out<=1;
   46011: out<=1;
   46012: out<=1;
   46013: out<=0;
   46014: out<=0;
   46015: out<=1;
   46016: out<=1;
   46017: out<=0;
   46018: out<=0;
   46019: out<=1;
   46020: out<=1;
   46021: out<=1;
   46022: out<=1;
   46023: out<=1;
   46024: out<=1;
   46025: out<=1;
   46026: out<=0;
   46027: out<=0;
   46028: out<=1;
   46029: out<=0;
   46030: out<=1;
   46031: out<=0;
   46032: out<=0;
   46033: out<=0;
   46034: out<=0;
   46035: out<=0;
   46036: out<=1;
   46037: out<=0;
   46038: out<=0;
   46039: out<=1;
   46040: out<=1;
   46041: out<=0;
   46042: out<=1;
   46043: out<=0;
   46044: out<=0;
   46045: out<=0;
   46046: out<=1;
   46047: out<=1;
   46048: out<=1;
   46049: out<=1;
   46050: out<=0;
   46051: out<=0;
   46052: out<=0;
   46053: out<=1;
   46054: out<=0;
   46055: out<=1;
   46056: out<=1;
   46057: out<=0;
   46058: out<=0;
   46059: out<=1;
   46060: out<=0;
   46061: out<=0;
   46062: out<=0;
   46063: out<=0;
   46064: out<=0;
   46065: out<=1;
   46066: out<=0;
   46067: out<=1;
   46068: out<=0;
   46069: out<=0;
   46070: out<=1;
   46071: out<=1;
   46072: out<=1;
   46073: out<=1;
   46074: out<=1;
   46075: out<=1;
   46076: out<=1;
   46077: out<=0;
   46078: out<=0;
   46079: out<=1;
   46080: out<=0;
   46081: out<=0;
   46082: out<=1;
   46083: out<=1;
   46084: out<=0;
   46085: out<=1;
   46086: out<=0;
   46087: out<=1;
   46088: out<=1;
   46089: out<=0;
   46090: out<=0;
   46091: out<=1;
   46092: out<=1;
   46093: out<=1;
   46094: out<=1;
   46095: out<=1;
   46096: out<=1;
   46097: out<=0;
   46098: out<=1;
   46099: out<=0;
   46100: out<=0;
   46101: out<=0;
   46102: out<=1;
   46103: out<=1;
   46104: out<=1;
   46105: out<=1;
   46106: out<=1;
   46107: out<=1;
   46108: out<=0;
   46109: out<=1;
   46110: out<=1;
   46111: out<=0;
   46112: out<=0;
   46113: out<=1;
   46114: out<=1;
   46115: out<=0;
   46116: out<=1;
   46117: out<=1;
   46118: out<=1;
   46119: out<=1;
   46120: out<=1;
   46121: out<=1;
   46122: out<=0;
   46123: out<=0;
   46124: out<=0;
   46125: out<=1;
   46126: out<=0;
   46127: out<=1;
   46128: out<=1;
   46129: out<=1;
   46130: out<=1;
   46131: out<=1;
   46132: out<=1;
   46133: out<=0;
   46134: out<=0;
   46135: out<=1;
   46136: out<=1;
   46137: out<=0;
   46138: out<=1;
   46139: out<=0;
   46140: out<=1;
   46141: out<=1;
   46142: out<=0;
   46143: out<=0;
   46144: out<=1;
   46145: out<=1;
   46146: out<=0;
   46147: out<=0;
   46148: out<=1;
   46149: out<=0;
   46150: out<=1;
   46151: out<=0;
   46152: out<=0;
   46153: out<=1;
   46154: out<=1;
   46155: out<=0;
   46156: out<=0;
   46157: out<=0;
   46158: out<=0;
   46159: out<=0;
   46160: out<=1;
   46161: out<=0;
   46162: out<=1;
   46163: out<=0;
   46164: out<=0;
   46165: out<=0;
   46166: out<=1;
   46167: out<=1;
   46168: out<=1;
   46169: out<=1;
   46170: out<=1;
   46171: out<=1;
   46172: out<=0;
   46173: out<=1;
   46174: out<=1;
   46175: out<=0;
   46176: out<=0;
   46177: out<=1;
   46178: out<=1;
   46179: out<=0;
   46180: out<=1;
   46181: out<=1;
   46182: out<=1;
   46183: out<=1;
   46184: out<=1;
   46185: out<=1;
   46186: out<=0;
   46187: out<=0;
   46188: out<=0;
   46189: out<=1;
   46190: out<=0;
   46191: out<=1;
   46192: out<=0;
   46193: out<=0;
   46194: out<=0;
   46195: out<=0;
   46196: out<=0;
   46197: out<=1;
   46198: out<=1;
   46199: out<=0;
   46200: out<=0;
   46201: out<=1;
   46202: out<=0;
   46203: out<=1;
   46204: out<=0;
   46205: out<=0;
   46206: out<=1;
   46207: out<=1;
   46208: out<=1;
   46209: out<=1;
   46210: out<=0;
   46211: out<=0;
   46212: out<=1;
   46213: out<=0;
   46214: out<=1;
   46215: out<=0;
   46216: out<=0;
   46217: out<=1;
   46218: out<=1;
   46219: out<=0;
   46220: out<=0;
   46221: out<=0;
   46222: out<=0;
   46223: out<=0;
   46224: out<=1;
   46225: out<=0;
   46226: out<=1;
   46227: out<=0;
   46228: out<=0;
   46229: out<=0;
   46230: out<=1;
   46231: out<=1;
   46232: out<=1;
   46233: out<=1;
   46234: out<=1;
   46235: out<=1;
   46236: out<=0;
   46237: out<=1;
   46238: out<=1;
   46239: out<=0;
   46240: out<=1;
   46241: out<=0;
   46242: out<=0;
   46243: out<=1;
   46244: out<=0;
   46245: out<=0;
   46246: out<=0;
   46247: out<=0;
   46248: out<=0;
   46249: out<=0;
   46250: out<=1;
   46251: out<=1;
   46252: out<=1;
   46253: out<=0;
   46254: out<=1;
   46255: out<=0;
   46256: out<=1;
   46257: out<=1;
   46258: out<=1;
   46259: out<=1;
   46260: out<=1;
   46261: out<=0;
   46262: out<=0;
   46263: out<=1;
   46264: out<=1;
   46265: out<=0;
   46266: out<=1;
   46267: out<=0;
   46268: out<=1;
   46269: out<=1;
   46270: out<=0;
   46271: out<=0;
   46272: out<=0;
   46273: out<=0;
   46274: out<=1;
   46275: out<=1;
   46276: out<=0;
   46277: out<=1;
   46278: out<=0;
   46279: out<=1;
   46280: out<=1;
   46281: out<=0;
   46282: out<=0;
   46283: out<=1;
   46284: out<=1;
   46285: out<=1;
   46286: out<=1;
   46287: out<=1;
   46288: out<=1;
   46289: out<=0;
   46290: out<=1;
   46291: out<=0;
   46292: out<=0;
   46293: out<=0;
   46294: out<=1;
   46295: out<=1;
   46296: out<=1;
   46297: out<=1;
   46298: out<=1;
   46299: out<=1;
   46300: out<=0;
   46301: out<=1;
   46302: out<=1;
   46303: out<=0;
   46304: out<=1;
   46305: out<=0;
   46306: out<=0;
   46307: out<=1;
   46308: out<=0;
   46309: out<=0;
   46310: out<=0;
   46311: out<=0;
   46312: out<=0;
   46313: out<=0;
   46314: out<=1;
   46315: out<=1;
   46316: out<=1;
   46317: out<=0;
   46318: out<=1;
   46319: out<=0;
   46320: out<=0;
   46321: out<=0;
   46322: out<=0;
   46323: out<=0;
   46324: out<=0;
   46325: out<=1;
   46326: out<=1;
   46327: out<=0;
   46328: out<=0;
   46329: out<=1;
   46330: out<=0;
   46331: out<=1;
   46332: out<=0;
   46333: out<=0;
   46334: out<=1;
   46335: out<=1;
   46336: out<=1;
   46337: out<=0;
   46338: out<=1;
   46339: out<=0;
   46340: out<=0;
   46341: out<=0;
   46342: out<=1;
   46343: out<=1;
   46344: out<=1;
   46345: out<=1;
   46346: out<=1;
   46347: out<=1;
   46348: out<=0;
   46349: out<=1;
   46350: out<=1;
   46351: out<=0;
   46352: out<=1;
   46353: out<=1;
   46354: out<=0;
   46355: out<=0;
   46356: out<=1;
   46357: out<=0;
   46358: out<=1;
   46359: out<=0;
   46360: out<=0;
   46361: out<=1;
   46362: out<=1;
   46363: out<=0;
   46364: out<=0;
   46365: out<=0;
   46366: out<=0;
   46367: out<=0;
   46368: out<=0;
   46369: out<=0;
   46370: out<=0;
   46371: out<=0;
   46372: out<=0;
   46373: out<=1;
   46374: out<=1;
   46375: out<=0;
   46376: out<=0;
   46377: out<=1;
   46378: out<=0;
   46379: out<=1;
   46380: out<=0;
   46381: out<=0;
   46382: out<=1;
   46383: out<=1;
   46384: out<=0;
   46385: out<=1;
   46386: out<=1;
   46387: out<=0;
   46388: out<=1;
   46389: out<=1;
   46390: out<=1;
   46391: out<=1;
   46392: out<=1;
   46393: out<=1;
   46394: out<=0;
   46395: out<=0;
   46396: out<=0;
   46397: out<=1;
   46398: out<=0;
   46399: out<=1;
   46400: out<=1;
   46401: out<=0;
   46402: out<=1;
   46403: out<=0;
   46404: out<=0;
   46405: out<=0;
   46406: out<=1;
   46407: out<=1;
   46408: out<=1;
   46409: out<=1;
   46410: out<=1;
   46411: out<=1;
   46412: out<=0;
   46413: out<=1;
   46414: out<=1;
   46415: out<=0;
   46416: out<=0;
   46417: out<=0;
   46418: out<=1;
   46419: out<=1;
   46420: out<=0;
   46421: out<=1;
   46422: out<=0;
   46423: out<=1;
   46424: out<=1;
   46425: out<=0;
   46426: out<=0;
   46427: out<=1;
   46428: out<=1;
   46429: out<=1;
   46430: out<=1;
   46431: out<=1;
   46432: out<=1;
   46433: out<=1;
   46434: out<=1;
   46435: out<=1;
   46436: out<=1;
   46437: out<=0;
   46438: out<=0;
   46439: out<=1;
   46440: out<=1;
   46441: out<=0;
   46442: out<=1;
   46443: out<=0;
   46444: out<=1;
   46445: out<=1;
   46446: out<=0;
   46447: out<=0;
   46448: out<=0;
   46449: out<=1;
   46450: out<=1;
   46451: out<=0;
   46452: out<=1;
   46453: out<=1;
   46454: out<=1;
   46455: out<=1;
   46456: out<=1;
   46457: out<=1;
   46458: out<=0;
   46459: out<=0;
   46460: out<=0;
   46461: out<=1;
   46462: out<=0;
   46463: out<=1;
   46464: out<=1;
   46465: out<=0;
   46466: out<=1;
   46467: out<=0;
   46468: out<=0;
   46469: out<=0;
   46470: out<=1;
   46471: out<=1;
   46472: out<=1;
   46473: out<=1;
   46474: out<=1;
   46475: out<=1;
   46476: out<=0;
   46477: out<=1;
   46478: out<=1;
   46479: out<=0;
   46480: out<=0;
   46481: out<=0;
   46482: out<=1;
   46483: out<=1;
   46484: out<=0;
   46485: out<=1;
   46486: out<=0;
   46487: out<=1;
   46488: out<=1;
   46489: out<=0;
   46490: out<=0;
   46491: out<=1;
   46492: out<=1;
   46493: out<=1;
   46494: out<=1;
   46495: out<=1;
   46496: out<=0;
   46497: out<=0;
   46498: out<=0;
   46499: out<=0;
   46500: out<=0;
   46501: out<=1;
   46502: out<=1;
   46503: out<=0;
   46504: out<=0;
   46505: out<=1;
   46506: out<=0;
   46507: out<=1;
   46508: out<=0;
   46509: out<=0;
   46510: out<=1;
   46511: out<=1;
   46512: out<=1;
   46513: out<=0;
   46514: out<=0;
   46515: out<=1;
   46516: out<=0;
   46517: out<=0;
   46518: out<=0;
   46519: out<=0;
   46520: out<=0;
   46521: out<=0;
   46522: out<=1;
   46523: out<=1;
   46524: out<=1;
   46525: out<=0;
   46526: out<=1;
   46527: out<=0;
   46528: out<=1;
   46529: out<=0;
   46530: out<=1;
   46531: out<=0;
   46532: out<=0;
   46533: out<=0;
   46534: out<=1;
   46535: out<=1;
   46536: out<=1;
   46537: out<=1;
   46538: out<=1;
   46539: out<=1;
   46540: out<=0;
   46541: out<=1;
   46542: out<=1;
   46543: out<=0;
   46544: out<=1;
   46545: out<=1;
   46546: out<=0;
   46547: out<=0;
   46548: out<=1;
   46549: out<=0;
   46550: out<=1;
   46551: out<=0;
   46552: out<=0;
   46553: out<=1;
   46554: out<=1;
   46555: out<=0;
   46556: out<=0;
   46557: out<=0;
   46558: out<=0;
   46559: out<=0;
   46560: out<=1;
   46561: out<=1;
   46562: out<=1;
   46563: out<=1;
   46564: out<=1;
   46565: out<=0;
   46566: out<=0;
   46567: out<=1;
   46568: out<=1;
   46569: out<=0;
   46570: out<=1;
   46571: out<=0;
   46572: out<=1;
   46573: out<=1;
   46574: out<=0;
   46575: out<=0;
   46576: out<=1;
   46577: out<=0;
   46578: out<=0;
   46579: out<=1;
   46580: out<=0;
   46581: out<=0;
   46582: out<=0;
   46583: out<=0;
   46584: out<=0;
   46585: out<=0;
   46586: out<=1;
   46587: out<=1;
   46588: out<=1;
   46589: out<=0;
   46590: out<=1;
   46591: out<=0;
   46592: out<=1;
   46593: out<=0;
   46594: out<=0;
   46595: out<=1;
   46596: out<=0;
   46597: out<=0;
   46598: out<=0;
   46599: out<=0;
   46600: out<=0;
   46601: out<=0;
   46602: out<=1;
   46603: out<=1;
   46604: out<=1;
   46605: out<=0;
   46606: out<=1;
   46607: out<=0;
   46608: out<=1;
   46609: out<=1;
   46610: out<=1;
   46611: out<=1;
   46612: out<=1;
   46613: out<=0;
   46614: out<=0;
   46615: out<=1;
   46616: out<=1;
   46617: out<=0;
   46618: out<=1;
   46619: out<=0;
   46620: out<=1;
   46621: out<=1;
   46622: out<=0;
   46623: out<=0;
   46624: out<=1;
   46625: out<=1;
   46626: out<=0;
   46627: out<=0;
   46628: out<=1;
   46629: out<=0;
   46630: out<=1;
   46631: out<=0;
   46632: out<=0;
   46633: out<=1;
   46634: out<=1;
   46635: out<=0;
   46636: out<=0;
   46637: out<=0;
   46638: out<=0;
   46639: out<=0;
   46640: out<=1;
   46641: out<=0;
   46642: out<=1;
   46643: out<=0;
   46644: out<=0;
   46645: out<=0;
   46646: out<=1;
   46647: out<=1;
   46648: out<=1;
   46649: out<=1;
   46650: out<=1;
   46651: out<=1;
   46652: out<=0;
   46653: out<=1;
   46654: out<=1;
   46655: out<=0;
   46656: out<=1;
   46657: out<=0;
   46658: out<=0;
   46659: out<=1;
   46660: out<=0;
   46661: out<=0;
   46662: out<=0;
   46663: out<=0;
   46664: out<=0;
   46665: out<=0;
   46666: out<=1;
   46667: out<=1;
   46668: out<=1;
   46669: out<=0;
   46670: out<=1;
   46671: out<=0;
   46672: out<=0;
   46673: out<=0;
   46674: out<=0;
   46675: out<=0;
   46676: out<=0;
   46677: out<=1;
   46678: out<=1;
   46679: out<=0;
   46680: out<=0;
   46681: out<=1;
   46682: out<=0;
   46683: out<=1;
   46684: out<=0;
   46685: out<=0;
   46686: out<=1;
   46687: out<=1;
   46688: out<=0;
   46689: out<=0;
   46690: out<=1;
   46691: out<=1;
   46692: out<=0;
   46693: out<=1;
   46694: out<=0;
   46695: out<=1;
   46696: out<=1;
   46697: out<=0;
   46698: out<=0;
   46699: out<=1;
   46700: out<=1;
   46701: out<=1;
   46702: out<=1;
   46703: out<=1;
   46704: out<=1;
   46705: out<=0;
   46706: out<=1;
   46707: out<=0;
   46708: out<=0;
   46709: out<=0;
   46710: out<=1;
   46711: out<=1;
   46712: out<=1;
   46713: out<=1;
   46714: out<=1;
   46715: out<=1;
   46716: out<=0;
   46717: out<=1;
   46718: out<=1;
   46719: out<=0;
   46720: out<=0;
   46721: out<=1;
   46722: out<=1;
   46723: out<=0;
   46724: out<=1;
   46725: out<=1;
   46726: out<=1;
   46727: out<=1;
   46728: out<=1;
   46729: out<=1;
   46730: out<=0;
   46731: out<=0;
   46732: out<=0;
   46733: out<=1;
   46734: out<=0;
   46735: out<=1;
   46736: out<=1;
   46737: out<=1;
   46738: out<=1;
   46739: out<=1;
   46740: out<=1;
   46741: out<=0;
   46742: out<=0;
   46743: out<=1;
   46744: out<=1;
   46745: out<=0;
   46746: out<=1;
   46747: out<=0;
   46748: out<=1;
   46749: out<=1;
   46750: out<=0;
   46751: out<=0;
   46752: out<=0;
   46753: out<=0;
   46754: out<=1;
   46755: out<=1;
   46756: out<=0;
   46757: out<=1;
   46758: out<=0;
   46759: out<=1;
   46760: out<=1;
   46761: out<=0;
   46762: out<=0;
   46763: out<=1;
   46764: out<=1;
   46765: out<=1;
   46766: out<=1;
   46767: out<=1;
   46768: out<=1;
   46769: out<=0;
   46770: out<=1;
   46771: out<=0;
   46772: out<=0;
   46773: out<=0;
   46774: out<=1;
   46775: out<=1;
   46776: out<=1;
   46777: out<=1;
   46778: out<=1;
   46779: out<=1;
   46780: out<=0;
   46781: out<=1;
   46782: out<=1;
   46783: out<=0;
   46784: out<=0;
   46785: out<=1;
   46786: out<=1;
   46787: out<=0;
   46788: out<=1;
   46789: out<=1;
   46790: out<=1;
   46791: out<=1;
   46792: out<=1;
   46793: out<=1;
   46794: out<=0;
   46795: out<=0;
   46796: out<=0;
   46797: out<=1;
   46798: out<=0;
   46799: out<=1;
   46800: out<=0;
   46801: out<=0;
   46802: out<=0;
   46803: out<=0;
   46804: out<=0;
   46805: out<=1;
   46806: out<=1;
   46807: out<=0;
   46808: out<=0;
   46809: out<=1;
   46810: out<=0;
   46811: out<=1;
   46812: out<=0;
   46813: out<=0;
   46814: out<=1;
   46815: out<=1;
   46816: out<=1;
   46817: out<=1;
   46818: out<=0;
   46819: out<=0;
   46820: out<=1;
   46821: out<=0;
   46822: out<=1;
   46823: out<=0;
   46824: out<=0;
   46825: out<=1;
   46826: out<=1;
   46827: out<=0;
   46828: out<=0;
   46829: out<=0;
   46830: out<=0;
   46831: out<=0;
   46832: out<=1;
   46833: out<=0;
   46834: out<=1;
   46835: out<=0;
   46836: out<=0;
   46837: out<=0;
   46838: out<=1;
   46839: out<=1;
   46840: out<=1;
   46841: out<=1;
   46842: out<=1;
   46843: out<=1;
   46844: out<=0;
   46845: out<=1;
   46846: out<=1;
   46847: out<=0;
   46848: out<=0;
   46849: out<=0;
   46850: out<=0;
   46851: out<=0;
   46852: out<=0;
   46853: out<=1;
   46854: out<=1;
   46855: out<=0;
   46856: out<=0;
   46857: out<=1;
   46858: out<=0;
   46859: out<=1;
   46860: out<=0;
   46861: out<=0;
   46862: out<=1;
   46863: out<=1;
   46864: out<=1;
   46865: out<=0;
   46866: out<=0;
   46867: out<=1;
   46868: out<=0;
   46869: out<=0;
   46870: out<=0;
   46871: out<=0;
   46872: out<=0;
   46873: out<=0;
   46874: out<=1;
   46875: out<=1;
   46876: out<=1;
   46877: out<=0;
   46878: out<=1;
   46879: out<=0;
   46880: out<=1;
   46881: out<=0;
   46882: out<=1;
   46883: out<=0;
   46884: out<=0;
   46885: out<=0;
   46886: out<=1;
   46887: out<=1;
   46888: out<=1;
   46889: out<=1;
   46890: out<=1;
   46891: out<=1;
   46892: out<=0;
   46893: out<=1;
   46894: out<=1;
   46895: out<=0;
   46896: out<=0;
   46897: out<=0;
   46898: out<=1;
   46899: out<=1;
   46900: out<=0;
   46901: out<=1;
   46902: out<=0;
   46903: out<=1;
   46904: out<=1;
   46905: out<=0;
   46906: out<=0;
   46907: out<=1;
   46908: out<=1;
   46909: out<=1;
   46910: out<=1;
   46911: out<=1;
   46912: out<=1;
   46913: out<=1;
   46914: out<=1;
   46915: out<=1;
   46916: out<=1;
   46917: out<=0;
   46918: out<=0;
   46919: out<=1;
   46920: out<=1;
   46921: out<=0;
   46922: out<=1;
   46923: out<=0;
   46924: out<=1;
   46925: out<=1;
   46926: out<=0;
   46927: out<=0;
   46928: out<=1;
   46929: out<=0;
   46930: out<=0;
   46931: out<=1;
   46932: out<=0;
   46933: out<=0;
   46934: out<=0;
   46935: out<=0;
   46936: out<=0;
   46937: out<=0;
   46938: out<=1;
   46939: out<=1;
   46940: out<=1;
   46941: out<=0;
   46942: out<=1;
   46943: out<=0;
   46944: out<=1;
   46945: out<=0;
   46946: out<=1;
   46947: out<=0;
   46948: out<=0;
   46949: out<=0;
   46950: out<=1;
   46951: out<=1;
   46952: out<=1;
   46953: out<=1;
   46954: out<=1;
   46955: out<=1;
   46956: out<=0;
   46957: out<=1;
   46958: out<=1;
   46959: out<=0;
   46960: out<=1;
   46961: out<=1;
   46962: out<=0;
   46963: out<=0;
   46964: out<=1;
   46965: out<=0;
   46966: out<=1;
   46967: out<=0;
   46968: out<=0;
   46969: out<=1;
   46970: out<=1;
   46971: out<=0;
   46972: out<=0;
   46973: out<=0;
   46974: out<=0;
   46975: out<=0;
   46976: out<=0;
   46977: out<=0;
   46978: out<=0;
   46979: out<=0;
   46980: out<=0;
   46981: out<=1;
   46982: out<=1;
   46983: out<=0;
   46984: out<=0;
   46985: out<=1;
   46986: out<=0;
   46987: out<=1;
   46988: out<=0;
   46989: out<=0;
   46990: out<=1;
   46991: out<=1;
   46992: out<=0;
   46993: out<=1;
   46994: out<=1;
   46995: out<=0;
   46996: out<=1;
   46997: out<=1;
   46998: out<=1;
   46999: out<=1;
   47000: out<=1;
   47001: out<=1;
   47002: out<=0;
   47003: out<=0;
   47004: out<=0;
   47005: out<=1;
   47006: out<=0;
   47007: out<=1;
   47008: out<=1;
   47009: out<=0;
   47010: out<=1;
   47011: out<=0;
   47012: out<=0;
   47013: out<=0;
   47014: out<=1;
   47015: out<=1;
   47016: out<=1;
   47017: out<=1;
   47018: out<=1;
   47019: out<=1;
   47020: out<=0;
   47021: out<=1;
   47022: out<=1;
   47023: out<=0;
   47024: out<=1;
   47025: out<=1;
   47026: out<=0;
   47027: out<=0;
   47028: out<=1;
   47029: out<=0;
   47030: out<=1;
   47031: out<=0;
   47032: out<=0;
   47033: out<=1;
   47034: out<=1;
   47035: out<=0;
   47036: out<=0;
   47037: out<=0;
   47038: out<=0;
   47039: out<=0;
   47040: out<=1;
   47041: out<=1;
   47042: out<=1;
   47043: out<=1;
   47044: out<=1;
   47045: out<=0;
   47046: out<=0;
   47047: out<=1;
   47048: out<=1;
   47049: out<=0;
   47050: out<=1;
   47051: out<=0;
   47052: out<=1;
   47053: out<=1;
   47054: out<=0;
   47055: out<=0;
   47056: out<=0;
   47057: out<=1;
   47058: out<=1;
   47059: out<=0;
   47060: out<=1;
   47061: out<=1;
   47062: out<=1;
   47063: out<=1;
   47064: out<=1;
   47065: out<=1;
   47066: out<=0;
   47067: out<=0;
   47068: out<=0;
   47069: out<=1;
   47070: out<=0;
   47071: out<=1;
   47072: out<=1;
   47073: out<=0;
   47074: out<=1;
   47075: out<=0;
   47076: out<=0;
   47077: out<=0;
   47078: out<=1;
   47079: out<=1;
   47080: out<=1;
   47081: out<=1;
   47082: out<=1;
   47083: out<=1;
   47084: out<=0;
   47085: out<=1;
   47086: out<=1;
   47087: out<=0;
   47088: out<=0;
   47089: out<=0;
   47090: out<=1;
   47091: out<=1;
   47092: out<=0;
   47093: out<=1;
   47094: out<=0;
   47095: out<=1;
   47096: out<=1;
   47097: out<=0;
   47098: out<=0;
   47099: out<=1;
   47100: out<=1;
   47101: out<=1;
   47102: out<=1;
   47103: out<=1;
   47104: out<=0;
   47105: out<=0;
   47106: out<=0;
   47107: out<=0;
   47108: out<=0;
   47109: out<=1;
   47110: out<=1;
   47111: out<=0;
   47112: out<=1;
   47113: out<=0;
   47114: out<=1;
   47115: out<=0;
   47116: out<=1;
   47117: out<=1;
   47118: out<=0;
   47119: out<=0;
   47120: out<=1;
   47121: out<=0;
   47122: out<=0;
   47123: out<=1;
   47124: out<=0;
   47125: out<=0;
   47126: out<=0;
   47127: out<=0;
   47128: out<=1;
   47129: out<=1;
   47130: out<=0;
   47131: out<=0;
   47132: out<=0;
   47133: out<=1;
   47134: out<=0;
   47135: out<=1;
   47136: out<=0;
   47137: out<=1;
   47138: out<=0;
   47139: out<=1;
   47140: out<=1;
   47141: out<=1;
   47142: out<=0;
   47143: out<=0;
   47144: out<=1;
   47145: out<=1;
   47146: out<=1;
   47147: out<=1;
   47148: out<=0;
   47149: out<=1;
   47150: out<=1;
   47151: out<=0;
   47152: out<=1;
   47153: out<=1;
   47154: out<=0;
   47155: out<=0;
   47156: out<=1;
   47157: out<=0;
   47158: out<=1;
   47159: out<=0;
   47160: out<=1;
   47161: out<=0;
   47162: out<=0;
   47163: out<=1;
   47164: out<=1;
   47165: out<=1;
   47166: out<=1;
   47167: out<=1;
   47168: out<=1;
   47169: out<=1;
   47170: out<=1;
   47171: out<=1;
   47172: out<=1;
   47173: out<=0;
   47174: out<=0;
   47175: out<=1;
   47176: out<=0;
   47177: out<=1;
   47178: out<=0;
   47179: out<=1;
   47180: out<=0;
   47181: out<=0;
   47182: out<=1;
   47183: out<=1;
   47184: out<=1;
   47185: out<=0;
   47186: out<=0;
   47187: out<=1;
   47188: out<=0;
   47189: out<=0;
   47190: out<=0;
   47191: out<=0;
   47192: out<=1;
   47193: out<=1;
   47194: out<=0;
   47195: out<=0;
   47196: out<=0;
   47197: out<=1;
   47198: out<=0;
   47199: out<=1;
   47200: out<=0;
   47201: out<=1;
   47202: out<=0;
   47203: out<=1;
   47204: out<=1;
   47205: out<=1;
   47206: out<=0;
   47207: out<=0;
   47208: out<=1;
   47209: out<=1;
   47210: out<=1;
   47211: out<=1;
   47212: out<=0;
   47213: out<=1;
   47214: out<=1;
   47215: out<=0;
   47216: out<=0;
   47217: out<=0;
   47218: out<=1;
   47219: out<=1;
   47220: out<=0;
   47221: out<=1;
   47222: out<=0;
   47223: out<=1;
   47224: out<=0;
   47225: out<=1;
   47226: out<=1;
   47227: out<=0;
   47228: out<=0;
   47229: out<=0;
   47230: out<=0;
   47231: out<=0;
   47232: out<=0;
   47233: out<=0;
   47234: out<=0;
   47235: out<=0;
   47236: out<=0;
   47237: out<=1;
   47238: out<=1;
   47239: out<=0;
   47240: out<=1;
   47241: out<=0;
   47242: out<=1;
   47243: out<=0;
   47244: out<=1;
   47245: out<=1;
   47246: out<=0;
   47247: out<=0;
   47248: out<=0;
   47249: out<=1;
   47250: out<=1;
   47251: out<=0;
   47252: out<=1;
   47253: out<=1;
   47254: out<=1;
   47255: out<=1;
   47256: out<=0;
   47257: out<=0;
   47258: out<=1;
   47259: out<=1;
   47260: out<=1;
   47261: out<=0;
   47262: out<=1;
   47263: out<=0;
   47264: out<=0;
   47265: out<=1;
   47266: out<=0;
   47267: out<=1;
   47268: out<=1;
   47269: out<=1;
   47270: out<=0;
   47271: out<=0;
   47272: out<=1;
   47273: out<=1;
   47274: out<=1;
   47275: out<=1;
   47276: out<=0;
   47277: out<=1;
   47278: out<=1;
   47279: out<=0;
   47280: out<=0;
   47281: out<=0;
   47282: out<=1;
   47283: out<=1;
   47284: out<=0;
   47285: out<=1;
   47286: out<=0;
   47287: out<=1;
   47288: out<=0;
   47289: out<=1;
   47290: out<=1;
   47291: out<=0;
   47292: out<=0;
   47293: out<=0;
   47294: out<=0;
   47295: out<=0;
   47296: out<=1;
   47297: out<=1;
   47298: out<=1;
   47299: out<=1;
   47300: out<=1;
   47301: out<=0;
   47302: out<=0;
   47303: out<=1;
   47304: out<=0;
   47305: out<=1;
   47306: out<=0;
   47307: out<=1;
   47308: out<=0;
   47309: out<=0;
   47310: out<=1;
   47311: out<=1;
   47312: out<=0;
   47313: out<=1;
   47314: out<=1;
   47315: out<=0;
   47316: out<=1;
   47317: out<=1;
   47318: out<=1;
   47319: out<=1;
   47320: out<=0;
   47321: out<=0;
   47322: out<=1;
   47323: out<=1;
   47324: out<=1;
   47325: out<=0;
   47326: out<=1;
   47327: out<=0;
   47328: out<=0;
   47329: out<=1;
   47330: out<=0;
   47331: out<=1;
   47332: out<=1;
   47333: out<=1;
   47334: out<=0;
   47335: out<=0;
   47336: out<=1;
   47337: out<=1;
   47338: out<=1;
   47339: out<=1;
   47340: out<=0;
   47341: out<=1;
   47342: out<=1;
   47343: out<=0;
   47344: out<=1;
   47345: out<=1;
   47346: out<=0;
   47347: out<=0;
   47348: out<=1;
   47349: out<=0;
   47350: out<=1;
   47351: out<=0;
   47352: out<=1;
   47353: out<=0;
   47354: out<=0;
   47355: out<=1;
   47356: out<=1;
   47357: out<=1;
   47358: out<=1;
   47359: out<=1;
   47360: out<=1;
   47361: out<=0;
   47362: out<=0;
   47363: out<=1;
   47364: out<=0;
   47365: out<=0;
   47366: out<=0;
   47367: out<=0;
   47368: out<=1;
   47369: out<=1;
   47370: out<=0;
   47371: out<=0;
   47372: out<=0;
   47373: out<=1;
   47374: out<=0;
   47375: out<=1;
   47376: out<=1;
   47377: out<=1;
   47378: out<=1;
   47379: out<=1;
   47380: out<=1;
   47381: out<=0;
   47382: out<=0;
   47383: out<=1;
   47384: out<=0;
   47385: out<=1;
   47386: out<=0;
   47387: out<=1;
   47388: out<=0;
   47389: out<=0;
   47390: out<=1;
   47391: out<=1;
   47392: out<=0;
   47393: out<=0;
   47394: out<=1;
   47395: out<=1;
   47396: out<=0;
   47397: out<=1;
   47398: out<=0;
   47399: out<=1;
   47400: out<=0;
   47401: out<=1;
   47402: out<=1;
   47403: out<=0;
   47404: out<=0;
   47405: out<=0;
   47406: out<=0;
   47407: out<=0;
   47408: out<=0;
   47409: out<=1;
   47410: out<=0;
   47411: out<=1;
   47412: out<=1;
   47413: out<=1;
   47414: out<=0;
   47415: out<=0;
   47416: out<=1;
   47417: out<=1;
   47418: out<=1;
   47419: out<=1;
   47420: out<=0;
   47421: out<=1;
   47422: out<=1;
   47423: out<=0;
   47424: out<=1;
   47425: out<=0;
   47426: out<=0;
   47427: out<=1;
   47428: out<=0;
   47429: out<=0;
   47430: out<=0;
   47431: out<=0;
   47432: out<=1;
   47433: out<=1;
   47434: out<=0;
   47435: out<=0;
   47436: out<=0;
   47437: out<=1;
   47438: out<=0;
   47439: out<=1;
   47440: out<=0;
   47441: out<=0;
   47442: out<=0;
   47443: out<=0;
   47444: out<=0;
   47445: out<=1;
   47446: out<=1;
   47447: out<=0;
   47448: out<=1;
   47449: out<=0;
   47450: out<=1;
   47451: out<=0;
   47452: out<=1;
   47453: out<=1;
   47454: out<=0;
   47455: out<=0;
   47456: out<=1;
   47457: out<=1;
   47458: out<=0;
   47459: out<=0;
   47460: out<=1;
   47461: out<=0;
   47462: out<=1;
   47463: out<=0;
   47464: out<=1;
   47465: out<=0;
   47466: out<=0;
   47467: out<=1;
   47468: out<=1;
   47469: out<=1;
   47470: out<=1;
   47471: out<=1;
   47472: out<=0;
   47473: out<=1;
   47474: out<=0;
   47475: out<=1;
   47476: out<=1;
   47477: out<=1;
   47478: out<=0;
   47479: out<=0;
   47480: out<=1;
   47481: out<=1;
   47482: out<=1;
   47483: out<=1;
   47484: out<=0;
   47485: out<=1;
   47486: out<=1;
   47487: out<=0;
   47488: out<=0;
   47489: out<=1;
   47490: out<=1;
   47491: out<=0;
   47492: out<=1;
   47493: out<=1;
   47494: out<=1;
   47495: out<=1;
   47496: out<=0;
   47497: out<=0;
   47498: out<=1;
   47499: out<=1;
   47500: out<=1;
   47501: out<=0;
   47502: out<=1;
   47503: out<=0;
   47504: out<=1;
   47505: out<=1;
   47506: out<=1;
   47507: out<=1;
   47508: out<=1;
   47509: out<=0;
   47510: out<=0;
   47511: out<=1;
   47512: out<=0;
   47513: out<=1;
   47514: out<=0;
   47515: out<=1;
   47516: out<=0;
   47517: out<=0;
   47518: out<=1;
   47519: out<=1;
   47520: out<=1;
   47521: out<=1;
   47522: out<=0;
   47523: out<=0;
   47524: out<=1;
   47525: out<=0;
   47526: out<=1;
   47527: out<=0;
   47528: out<=1;
   47529: out<=0;
   47530: out<=0;
   47531: out<=1;
   47532: out<=1;
   47533: out<=1;
   47534: out<=1;
   47535: out<=1;
   47536: out<=0;
   47537: out<=1;
   47538: out<=0;
   47539: out<=1;
   47540: out<=1;
   47541: out<=1;
   47542: out<=0;
   47543: out<=0;
   47544: out<=1;
   47545: out<=1;
   47546: out<=1;
   47547: out<=1;
   47548: out<=0;
   47549: out<=1;
   47550: out<=1;
   47551: out<=0;
   47552: out<=0;
   47553: out<=1;
   47554: out<=1;
   47555: out<=0;
   47556: out<=1;
   47557: out<=1;
   47558: out<=1;
   47559: out<=1;
   47560: out<=0;
   47561: out<=0;
   47562: out<=1;
   47563: out<=1;
   47564: out<=1;
   47565: out<=0;
   47566: out<=1;
   47567: out<=0;
   47568: out<=0;
   47569: out<=0;
   47570: out<=0;
   47571: out<=0;
   47572: out<=0;
   47573: out<=1;
   47574: out<=1;
   47575: out<=0;
   47576: out<=1;
   47577: out<=0;
   47578: out<=1;
   47579: out<=0;
   47580: out<=1;
   47581: out<=1;
   47582: out<=0;
   47583: out<=0;
   47584: out<=0;
   47585: out<=0;
   47586: out<=1;
   47587: out<=1;
   47588: out<=0;
   47589: out<=1;
   47590: out<=0;
   47591: out<=1;
   47592: out<=0;
   47593: out<=1;
   47594: out<=1;
   47595: out<=0;
   47596: out<=0;
   47597: out<=0;
   47598: out<=0;
   47599: out<=0;
   47600: out<=0;
   47601: out<=1;
   47602: out<=0;
   47603: out<=1;
   47604: out<=1;
   47605: out<=1;
   47606: out<=0;
   47607: out<=0;
   47608: out<=1;
   47609: out<=1;
   47610: out<=1;
   47611: out<=1;
   47612: out<=0;
   47613: out<=1;
   47614: out<=1;
   47615: out<=0;
   47616: out<=0;
   47617: out<=1;
   47618: out<=0;
   47619: out<=1;
   47620: out<=1;
   47621: out<=1;
   47622: out<=0;
   47623: out<=0;
   47624: out<=1;
   47625: out<=1;
   47626: out<=1;
   47627: out<=1;
   47628: out<=0;
   47629: out<=1;
   47630: out<=1;
   47631: out<=0;
   47632: out<=0;
   47633: out<=0;
   47634: out<=1;
   47635: out<=1;
   47636: out<=0;
   47637: out<=1;
   47638: out<=0;
   47639: out<=1;
   47640: out<=0;
   47641: out<=1;
   47642: out<=1;
   47643: out<=0;
   47644: out<=0;
   47645: out<=0;
   47646: out<=0;
   47647: out<=0;
   47648: out<=0;
   47649: out<=0;
   47650: out<=0;
   47651: out<=0;
   47652: out<=0;
   47653: out<=1;
   47654: out<=1;
   47655: out<=0;
   47656: out<=1;
   47657: out<=0;
   47658: out<=1;
   47659: out<=0;
   47660: out<=1;
   47661: out<=1;
   47662: out<=0;
   47663: out<=0;
   47664: out<=0;
   47665: out<=1;
   47666: out<=1;
   47667: out<=0;
   47668: out<=1;
   47669: out<=1;
   47670: out<=1;
   47671: out<=1;
   47672: out<=0;
   47673: out<=0;
   47674: out<=1;
   47675: out<=1;
   47676: out<=1;
   47677: out<=0;
   47678: out<=1;
   47679: out<=0;
   47680: out<=0;
   47681: out<=1;
   47682: out<=0;
   47683: out<=1;
   47684: out<=1;
   47685: out<=1;
   47686: out<=0;
   47687: out<=0;
   47688: out<=1;
   47689: out<=1;
   47690: out<=1;
   47691: out<=1;
   47692: out<=0;
   47693: out<=1;
   47694: out<=1;
   47695: out<=0;
   47696: out<=1;
   47697: out<=1;
   47698: out<=0;
   47699: out<=0;
   47700: out<=1;
   47701: out<=0;
   47702: out<=1;
   47703: out<=0;
   47704: out<=1;
   47705: out<=0;
   47706: out<=0;
   47707: out<=1;
   47708: out<=1;
   47709: out<=1;
   47710: out<=1;
   47711: out<=1;
   47712: out<=1;
   47713: out<=1;
   47714: out<=1;
   47715: out<=1;
   47716: out<=1;
   47717: out<=0;
   47718: out<=0;
   47719: out<=1;
   47720: out<=0;
   47721: out<=1;
   47722: out<=0;
   47723: out<=1;
   47724: out<=0;
   47725: out<=0;
   47726: out<=1;
   47727: out<=1;
   47728: out<=0;
   47729: out<=1;
   47730: out<=1;
   47731: out<=0;
   47732: out<=1;
   47733: out<=1;
   47734: out<=1;
   47735: out<=1;
   47736: out<=0;
   47737: out<=0;
   47738: out<=1;
   47739: out<=1;
   47740: out<=1;
   47741: out<=0;
   47742: out<=1;
   47743: out<=0;
   47744: out<=0;
   47745: out<=1;
   47746: out<=0;
   47747: out<=1;
   47748: out<=1;
   47749: out<=1;
   47750: out<=0;
   47751: out<=0;
   47752: out<=1;
   47753: out<=1;
   47754: out<=1;
   47755: out<=1;
   47756: out<=0;
   47757: out<=1;
   47758: out<=1;
   47759: out<=0;
   47760: out<=1;
   47761: out<=1;
   47762: out<=0;
   47763: out<=0;
   47764: out<=1;
   47765: out<=0;
   47766: out<=1;
   47767: out<=0;
   47768: out<=1;
   47769: out<=0;
   47770: out<=0;
   47771: out<=1;
   47772: out<=1;
   47773: out<=1;
   47774: out<=1;
   47775: out<=1;
   47776: out<=0;
   47777: out<=0;
   47778: out<=0;
   47779: out<=0;
   47780: out<=0;
   47781: out<=1;
   47782: out<=1;
   47783: out<=0;
   47784: out<=1;
   47785: out<=0;
   47786: out<=1;
   47787: out<=0;
   47788: out<=1;
   47789: out<=1;
   47790: out<=0;
   47791: out<=0;
   47792: out<=1;
   47793: out<=0;
   47794: out<=0;
   47795: out<=1;
   47796: out<=0;
   47797: out<=0;
   47798: out<=0;
   47799: out<=0;
   47800: out<=1;
   47801: out<=1;
   47802: out<=0;
   47803: out<=0;
   47804: out<=0;
   47805: out<=1;
   47806: out<=0;
   47807: out<=1;
   47808: out<=0;
   47809: out<=1;
   47810: out<=0;
   47811: out<=1;
   47812: out<=1;
   47813: out<=1;
   47814: out<=0;
   47815: out<=0;
   47816: out<=1;
   47817: out<=1;
   47818: out<=1;
   47819: out<=1;
   47820: out<=0;
   47821: out<=1;
   47822: out<=1;
   47823: out<=0;
   47824: out<=0;
   47825: out<=0;
   47826: out<=1;
   47827: out<=1;
   47828: out<=0;
   47829: out<=1;
   47830: out<=0;
   47831: out<=1;
   47832: out<=0;
   47833: out<=1;
   47834: out<=1;
   47835: out<=0;
   47836: out<=0;
   47837: out<=0;
   47838: out<=0;
   47839: out<=0;
   47840: out<=1;
   47841: out<=1;
   47842: out<=1;
   47843: out<=1;
   47844: out<=1;
   47845: out<=0;
   47846: out<=0;
   47847: out<=1;
   47848: out<=0;
   47849: out<=1;
   47850: out<=0;
   47851: out<=1;
   47852: out<=0;
   47853: out<=0;
   47854: out<=1;
   47855: out<=1;
   47856: out<=1;
   47857: out<=0;
   47858: out<=0;
   47859: out<=1;
   47860: out<=0;
   47861: out<=0;
   47862: out<=0;
   47863: out<=0;
   47864: out<=1;
   47865: out<=1;
   47866: out<=0;
   47867: out<=0;
   47868: out<=0;
   47869: out<=1;
   47870: out<=0;
   47871: out<=1;
   47872: out<=1;
   47873: out<=1;
   47874: out<=0;
   47875: out<=0;
   47876: out<=1;
   47877: out<=0;
   47878: out<=1;
   47879: out<=0;
   47880: out<=1;
   47881: out<=0;
   47882: out<=0;
   47883: out<=1;
   47884: out<=1;
   47885: out<=1;
   47886: out<=1;
   47887: out<=1;
   47888: out<=0;
   47889: out<=1;
   47890: out<=0;
   47891: out<=1;
   47892: out<=1;
   47893: out<=1;
   47894: out<=0;
   47895: out<=0;
   47896: out<=1;
   47897: out<=1;
   47898: out<=1;
   47899: out<=1;
   47900: out<=0;
   47901: out<=1;
   47902: out<=1;
   47903: out<=0;
   47904: out<=0;
   47905: out<=1;
   47906: out<=1;
   47907: out<=0;
   47908: out<=1;
   47909: out<=1;
   47910: out<=1;
   47911: out<=1;
   47912: out<=0;
   47913: out<=0;
   47914: out<=1;
   47915: out<=1;
   47916: out<=1;
   47917: out<=0;
   47918: out<=1;
   47919: out<=0;
   47920: out<=1;
   47921: out<=1;
   47922: out<=1;
   47923: out<=1;
   47924: out<=1;
   47925: out<=0;
   47926: out<=0;
   47927: out<=1;
   47928: out<=0;
   47929: out<=1;
   47930: out<=0;
   47931: out<=1;
   47932: out<=0;
   47933: out<=0;
   47934: out<=1;
   47935: out<=1;
   47936: out<=0;
   47937: out<=0;
   47938: out<=1;
   47939: out<=1;
   47940: out<=0;
   47941: out<=1;
   47942: out<=0;
   47943: out<=1;
   47944: out<=0;
   47945: out<=1;
   47946: out<=1;
   47947: out<=0;
   47948: out<=0;
   47949: out<=0;
   47950: out<=0;
   47951: out<=0;
   47952: out<=0;
   47953: out<=1;
   47954: out<=0;
   47955: out<=1;
   47956: out<=1;
   47957: out<=1;
   47958: out<=0;
   47959: out<=0;
   47960: out<=1;
   47961: out<=1;
   47962: out<=1;
   47963: out<=1;
   47964: out<=0;
   47965: out<=1;
   47966: out<=1;
   47967: out<=0;
   47968: out<=0;
   47969: out<=1;
   47970: out<=1;
   47971: out<=0;
   47972: out<=1;
   47973: out<=1;
   47974: out<=1;
   47975: out<=1;
   47976: out<=0;
   47977: out<=0;
   47978: out<=1;
   47979: out<=1;
   47980: out<=1;
   47981: out<=0;
   47982: out<=1;
   47983: out<=0;
   47984: out<=0;
   47985: out<=0;
   47986: out<=0;
   47987: out<=0;
   47988: out<=0;
   47989: out<=1;
   47990: out<=1;
   47991: out<=0;
   47992: out<=1;
   47993: out<=0;
   47994: out<=1;
   47995: out<=0;
   47996: out<=1;
   47997: out<=1;
   47998: out<=0;
   47999: out<=0;
   48000: out<=0;
   48001: out<=0;
   48002: out<=1;
   48003: out<=1;
   48004: out<=0;
   48005: out<=1;
   48006: out<=0;
   48007: out<=1;
   48008: out<=0;
   48009: out<=1;
   48010: out<=1;
   48011: out<=0;
   48012: out<=0;
   48013: out<=0;
   48014: out<=0;
   48015: out<=0;
   48016: out<=0;
   48017: out<=1;
   48018: out<=0;
   48019: out<=1;
   48020: out<=1;
   48021: out<=1;
   48022: out<=0;
   48023: out<=0;
   48024: out<=1;
   48025: out<=1;
   48026: out<=1;
   48027: out<=1;
   48028: out<=0;
   48029: out<=1;
   48030: out<=1;
   48031: out<=0;
   48032: out<=1;
   48033: out<=0;
   48034: out<=0;
   48035: out<=1;
   48036: out<=0;
   48037: out<=0;
   48038: out<=0;
   48039: out<=0;
   48040: out<=1;
   48041: out<=1;
   48042: out<=0;
   48043: out<=0;
   48044: out<=0;
   48045: out<=1;
   48046: out<=0;
   48047: out<=1;
   48048: out<=1;
   48049: out<=1;
   48050: out<=1;
   48051: out<=1;
   48052: out<=1;
   48053: out<=0;
   48054: out<=0;
   48055: out<=1;
   48056: out<=0;
   48057: out<=1;
   48058: out<=0;
   48059: out<=1;
   48060: out<=0;
   48061: out<=0;
   48062: out<=1;
   48063: out<=1;
   48064: out<=1;
   48065: out<=1;
   48066: out<=0;
   48067: out<=0;
   48068: out<=1;
   48069: out<=0;
   48070: out<=1;
   48071: out<=0;
   48072: out<=1;
   48073: out<=0;
   48074: out<=0;
   48075: out<=1;
   48076: out<=1;
   48077: out<=1;
   48078: out<=1;
   48079: out<=1;
   48080: out<=0;
   48081: out<=1;
   48082: out<=0;
   48083: out<=1;
   48084: out<=1;
   48085: out<=1;
   48086: out<=0;
   48087: out<=0;
   48088: out<=1;
   48089: out<=1;
   48090: out<=1;
   48091: out<=1;
   48092: out<=0;
   48093: out<=1;
   48094: out<=1;
   48095: out<=0;
   48096: out<=1;
   48097: out<=0;
   48098: out<=0;
   48099: out<=1;
   48100: out<=0;
   48101: out<=0;
   48102: out<=0;
   48103: out<=0;
   48104: out<=1;
   48105: out<=1;
   48106: out<=0;
   48107: out<=0;
   48108: out<=0;
   48109: out<=1;
   48110: out<=0;
   48111: out<=1;
   48112: out<=0;
   48113: out<=0;
   48114: out<=0;
   48115: out<=0;
   48116: out<=0;
   48117: out<=1;
   48118: out<=1;
   48119: out<=0;
   48120: out<=1;
   48121: out<=0;
   48122: out<=1;
   48123: out<=0;
   48124: out<=1;
   48125: out<=1;
   48126: out<=0;
   48127: out<=0;
   48128: out<=0;
   48129: out<=1;
   48130: out<=1;
   48131: out<=0;
   48132: out<=0;
   48133: out<=0;
   48134: out<=0;
   48135: out<=0;
   48136: out<=1;
   48137: out<=1;
   48138: out<=0;
   48139: out<=0;
   48140: out<=1;
   48141: out<=0;
   48142: out<=1;
   48143: out<=0;
   48144: out<=1;
   48145: out<=1;
   48146: out<=1;
   48147: out<=1;
   48148: out<=0;
   48149: out<=1;
   48150: out<=1;
   48151: out<=0;
   48152: out<=1;
   48153: out<=0;
   48154: out<=1;
   48155: out<=0;
   48156: out<=0;
   48157: out<=0;
   48158: out<=1;
   48159: out<=1;
   48160: out<=0;
   48161: out<=0;
   48162: out<=1;
   48163: out<=1;
   48164: out<=1;
   48165: out<=0;
   48166: out<=1;
   48167: out<=0;
   48168: out<=1;
   48169: out<=0;
   48170: out<=0;
   48171: out<=1;
   48172: out<=0;
   48173: out<=0;
   48174: out<=0;
   48175: out<=0;
   48176: out<=1;
   48177: out<=0;
   48178: out<=1;
   48179: out<=0;
   48180: out<=1;
   48181: out<=1;
   48182: out<=0;
   48183: out<=0;
   48184: out<=1;
   48185: out<=1;
   48186: out<=1;
   48187: out<=1;
   48188: out<=1;
   48189: out<=0;
   48190: out<=0;
   48191: out<=1;
   48192: out<=0;
   48193: out<=1;
   48194: out<=1;
   48195: out<=0;
   48196: out<=0;
   48197: out<=0;
   48198: out<=0;
   48199: out<=0;
   48200: out<=1;
   48201: out<=1;
   48202: out<=0;
   48203: out<=0;
   48204: out<=1;
   48205: out<=0;
   48206: out<=1;
   48207: out<=0;
   48208: out<=0;
   48209: out<=0;
   48210: out<=0;
   48211: out<=0;
   48212: out<=1;
   48213: out<=0;
   48214: out<=0;
   48215: out<=1;
   48216: out<=0;
   48217: out<=1;
   48218: out<=0;
   48219: out<=1;
   48220: out<=1;
   48221: out<=1;
   48222: out<=0;
   48223: out<=0;
   48224: out<=1;
   48225: out<=1;
   48226: out<=0;
   48227: out<=0;
   48228: out<=0;
   48229: out<=1;
   48230: out<=0;
   48231: out<=1;
   48232: out<=0;
   48233: out<=1;
   48234: out<=1;
   48235: out<=0;
   48236: out<=1;
   48237: out<=1;
   48238: out<=1;
   48239: out<=1;
   48240: out<=1;
   48241: out<=0;
   48242: out<=1;
   48243: out<=0;
   48244: out<=1;
   48245: out<=1;
   48246: out<=0;
   48247: out<=0;
   48248: out<=1;
   48249: out<=1;
   48250: out<=1;
   48251: out<=1;
   48252: out<=1;
   48253: out<=0;
   48254: out<=0;
   48255: out<=1;
   48256: out<=1;
   48257: out<=0;
   48258: out<=0;
   48259: out<=1;
   48260: out<=1;
   48261: out<=1;
   48262: out<=1;
   48263: out<=1;
   48264: out<=0;
   48265: out<=0;
   48266: out<=1;
   48267: out<=1;
   48268: out<=0;
   48269: out<=1;
   48270: out<=0;
   48271: out<=1;
   48272: out<=1;
   48273: out<=1;
   48274: out<=1;
   48275: out<=1;
   48276: out<=0;
   48277: out<=1;
   48278: out<=1;
   48279: out<=0;
   48280: out<=1;
   48281: out<=0;
   48282: out<=1;
   48283: out<=0;
   48284: out<=0;
   48285: out<=0;
   48286: out<=1;
   48287: out<=1;
   48288: out<=1;
   48289: out<=1;
   48290: out<=0;
   48291: out<=0;
   48292: out<=0;
   48293: out<=1;
   48294: out<=0;
   48295: out<=1;
   48296: out<=0;
   48297: out<=1;
   48298: out<=1;
   48299: out<=0;
   48300: out<=1;
   48301: out<=1;
   48302: out<=1;
   48303: out<=1;
   48304: out<=1;
   48305: out<=0;
   48306: out<=1;
   48307: out<=0;
   48308: out<=1;
   48309: out<=1;
   48310: out<=0;
   48311: out<=0;
   48312: out<=1;
   48313: out<=1;
   48314: out<=1;
   48315: out<=1;
   48316: out<=1;
   48317: out<=0;
   48318: out<=0;
   48319: out<=1;
   48320: out<=1;
   48321: out<=0;
   48322: out<=0;
   48323: out<=1;
   48324: out<=1;
   48325: out<=1;
   48326: out<=1;
   48327: out<=1;
   48328: out<=0;
   48329: out<=0;
   48330: out<=1;
   48331: out<=1;
   48332: out<=0;
   48333: out<=1;
   48334: out<=0;
   48335: out<=1;
   48336: out<=0;
   48337: out<=0;
   48338: out<=0;
   48339: out<=0;
   48340: out<=1;
   48341: out<=0;
   48342: out<=0;
   48343: out<=1;
   48344: out<=0;
   48345: out<=1;
   48346: out<=0;
   48347: out<=1;
   48348: out<=1;
   48349: out<=1;
   48350: out<=0;
   48351: out<=0;
   48352: out<=0;
   48353: out<=0;
   48354: out<=1;
   48355: out<=1;
   48356: out<=1;
   48357: out<=0;
   48358: out<=1;
   48359: out<=0;
   48360: out<=1;
   48361: out<=0;
   48362: out<=0;
   48363: out<=1;
   48364: out<=0;
   48365: out<=0;
   48366: out<=0;
   48367: out<=0;
   48368: out<=1;
   48369: out<=0;
   48370: out<=1;
   48371: out<=0;
   48372: out<=1;
   48373: out<=1;
   48374: out<=0;
   48375: out<=0;
   48376: out<=1;
   48377: out<=1;
   48378: out<=1;
   48379: out<=1;
   48380: out<=1;
   48381: out<=0;
   48382: out<=0;
   48383: out<=1;
   48384: out<=0;
   48385: out<=0;
   48386: out<=0;
   48387: out<=0;
   48388: out<=1;
   48389: out<=0;
   48390: out<=0;
   48391: out<=1;
   48392: out<=0;
   48393: out<=1;
   48394: out<=0;
   48395: out<=1;
   48396: out<=1;
   48397: out<=1;
   48398: out<=0;
   48399: out<=0;
   48400: out<=0;
   48401: out<=1;
   48402: out<=1;
   48403: out<=0;
   48404: out<=0;
   48405: out<=0;
   48406: out<=0;
   48407: out<=0;
   48408: out<=1;
   48409: out<=1;
   48410: out<=0;
   48411: out<=0;
   48412: out<=1;
   48413: out<=0;
   48414: out<=1;
   48415: out<=0;
   48416: out<=1;
   48417: out<=0;
   48418: out<=1;
   48419: out<=0;
   48420: out<=1;
   48421: out<=1;
   48422: out<=0;
   48423: out<=0;
   48424: out<=1;
   48425: out<=1;
   48426: out<=1;
   48427: out<=1;
   48428: out<=1;
   48429: out<=0;
   48430: out<=0;
   48431: out<=1;
   48432: out<=1;
   48433: out<=1;
   48434: out<=0;
   48435: out<=0;
   48436: out<=0;
   48437: out<=1;
   48438: out<=0;
   48439: out<=1;
   48440: out<=0;
   48441: out<=1;
   48442: out<=1;
   48443: out<=0;
   48444: out<=1;
   48445: out<=1;
   48446: out<=1;
   48447: out<=1;
   48448: out<=1;
   48449: out<=1;
   48450: out<=1;
   48451: out<=1;
   48452: out<=0;
   48453: out<=1;
   48454: out<=1;
   48455: out<=0;
   48456: out<=1;
   48457: out<=0;
   48458: out<=1;
   48459: out<=0;
   48460: out<=0;
   48461: out<=0;
   48462: out<=1;
   48463: out<=1;
   48464: out<=0;
   48465: out<=1;
   48466: out<=1;
   48467: out<=0;
   48468: out<=0;
   48469: out<=0;
   48470: out<=0;
   48471: out<=0;
   48472: out<=1;
   48473: out<=1;
   48474: out<=0;
   48475: out<=0;
   48476: out<=1;
   48477: out<=0;
   48478: out<=1;
   48479: out<=0;
   48480: out<=1;
   48481: out<=0;
   48482: out<=1;
   48483: out<=0;
   48484: out<=1;
   48485: out<=1;
   48486: out<=0;
   48487: out<=0;
   48488: out<=1;
   48489: out<=1;
   48490: out<=1;
   48491: out<=1;
   48492: out<=1;
   48493: out<=0;
   48494: out<=0;
   48495: out<=1;
   48496: out<=0;
   48497: out<=0;
   48498: out<=1;
   48499: out<=1;
   48500: out<=1;
   48501: out<=0;
   48502: out<=1;
   48503: out<=0;
   48504: out<=1;
   48505: out<=0;
   48506: out<=0;
   48507: out<=1;
   48508: out<=0;
   48509: out<=0;
   48510: out<=0;
   48511: out<=0;
   48512: out<=0;
   48513: out<=0;
   48514: out<=0;
   48515: out<=0;
   48516: out<=1;
   48517: out<=0;
   48518: out<=0;
   48519: out<=1;
   48520: out<=0;
   48521: out<=1;
   48522: out<=0;
   48523: out<=1;
   48524: out<=1;
   48525: out<=1;
   48526: out<=0;
   48527: out<=0;
   48528: out<=1;
   48529: out<=0;
   48530: out<=0;
   48531: out<=1;
   48532: out<=1;
   48533: out<=1;
   48534: out<=1;
   48535: out<=1;
   48536: out<=0;
   48537: out<=0;
   48538: out<=1;
   48539: out<=1;
   48540: out<=0;
   48541: out<=1;
   48542: out<=0;
   48543: out<=1;
   48544: out<=1;
   48545: out<=0;
   48546: out<=1;
   48547: out<=0;
   48548: out<=1;
   48549: out<=1;
   48550: out<=0;
   48551: out<=0;
   48552: out<=1;
   48553: out<=1;
   48554: out<=1;
   48555: out<=1;
   48556: out<=1;
   48557: out<=0;
   48558: out<=0;
   48559: out<=1;
   48560: out<=0;
   48561: out<=0;
   48562: out<=1;
   48563: out<=1;
   48564: out<=1;
   48565: out<=0;
   48566: out<=1;
   48567: out<=0;
   48568: out<=1;
   48569: out<=0;
   48570: out<=0;
   48571: out<=1;
   48572: out<=0;
   48573: out<=0;
   48574: out<=0;
   48575: out<=0;
   48576: out<=1;
   48577: out<=1;
   48578: out<=1;
   48579: out<=1;
   48580: out<=0;
   48581: out<=1;
   48582: out<=1;
   48583: out<=0;
   48584: out<=1;
   48585: out<=0;
   48586: out<=1;
   48587: out<=0;
   48588: out<=0;
   48589: out<=0;
   48590: out<=1;
   48591: out<=1;
   48592: out<=1;
   48593: out<=0;
   48594: out<=0;
   48595: out<=1;
   48596: out<=1;
   48597: out<=1;
   48598: out<=1;
   48599: out<=1;
   48600: out<=0;
   48601: out<=0;
   48602: out<=1;
   48603: out<=1;
   48604: out<=0;
   48605: out<=1;
   48606: out<=0;
   48607: out<=1;
   48608: out<=1;
   48609: out<=0;
   48610: out<=1;
   48611: out<=0;
   48612: out<=1;
   48613: out<=1;
   48614: out<=0;
   48615: out<=0;
   48616: out<=1;
   48617: out<=1;
   48618: out<=1;
   48619: out<=1;
   48620: out<=1;
   48621: out<=0;
   48622: out<=0;
   48623: out<=1;
   48624: out<=1;
   48625: out<=1;
   48626: out<=0;
   48627: out<=0;
   48628: out<=0;
   48629: out<=1;
   48630: out<=0;
   48631: out<=1;
   48632: out<=0;
   48633: out<=1;
   48634: out<=1;
   48635: out<=0;
   48636: out<=1;
   48637: out<=1;
   48638: out<=1;
   48639: out<=1;
   48640: out<=1;
   48641: out<=1;
   48642: out<=0;
   48643: out<=0;
   48644: out<=0;
   48645: out<=1;
   48646: out<=0;
   48647: out<=1;
   48648: out<=0;
   48649: out<=1;
   48650: out<=1;
   48651: out<=0;
   48652: out<=1;
   48653: out<=1;
   48654: out<=1;
   48655: out<=1;
   48656: out<=1;
   48657: out<=0;
   48658: out<=1;
   48659: out<=0;
   48660: out<=1;
   48661: out<=1;
   48662: out<=0;
   48663: out<=0;
   48664: out<=1;
   48665: out<=1;
   48666: out<=1;
   48667: out<=1;
   48668: out<=1;
   48669: out<=0;
   48670: out<=0;
   48671: out<=1;
   48672: out<=1;
   48673: out<=0;
   48674: out<=0;
   48675: out<=1;
   48676: out<=1;
   48677: out<=1;
   48678: out<=1;
   48679: out<=1;
   48680: out<=0;
   48681: out<=0;
   48682: out<=1;
   48683: out<=1;
   48684: out<=0;
   48685: out<=1;
   48686: out<=0;
   48687: out<=1;
   48688: out<=1;
   48689: out<=1;
   48690: out<=1;
   48691: out<=1;
   48692: out<=0;
   48693: out<=1;
   48694: out<=1;
   48695: out<=0;
   48696: out<=1;
   48697: out<=0;
   48698: out<=1;
   48699: out<=0;
   48700: out<=0;
   48701: out<=0;
   48702: out<=1;
   48703: out<=1;
   48704: out<=0;
   48705: out<=0;
   48706: out<=1;
   48707: out<=1;
   48708: out<=1;
   48709: out<=0;
   48710: out<=1;
   48711: out<=0;
   48712: out<=1;
   48713: out<=0;
   48714: out<=0;
   48715: out<=1;
   48716: out<=0;
   48717: out<=0;
   48718: out<=0;
   48719: out<=0;
   48720: out<=1;
   48721: out<=0;
   48722: out<=1;
   48723: out<=0;
   48724: out<=1;
   48725: out<=1;
   48726: out<=0;
   48727: out<=0;
   48728: out<=1;
   48729: out<=1;
   48730: out<=1;
   48731: out<=1;
   48732: out<=1;
   48733: out<=0;
   48734: out<=0;
   48735: out<=1;
   48736: out<=1;
   48737: out<=0;
   48738: out<=0;
   48739: out<=1;
   48740: out<=1;
   48741: out<=1;
   48742: out<=1;
   48743: out<=1;
   48744: out<=0;
   48745: out<=0;
   48746: out<=1;
   48747: out<=1;
   48748: out<=0;
   48749: out<=1;
   48750: out<=0;
   48751: out<=1;
   48752: out<=0;
   48753: out<=0;
   48754: out<=0;
   48755: out<=0;
   48756: out<=1;
   48757: out<=0;
   48758: out<=0;
   48759: out<=1;
   48760: out<=0;
   48761: out<=1;
   48762: out<=0;
   48763: out<=1;
   48764: out<=1;
   48765: out<=1;
   48766: out<=0;
   48767: out<=0;
   48768: out<=0;
   48769: out<=0;
   48770: out<=1;
   48771: out<=1;
   48772: out<=1;
   48773: out<=0;
   48774: out<=1;
   48775: out<=0;
   48776: out<=1;
   48777: out<=0;
   48778: out<=0;
   48779: out<=1;
   48780: out<=0;
   48781: out<=0;
   48782: out<=0;
   48783: out<=0;
   48784: out<=1;
   48785: out<=0;
   48786: out<=1;
   48787: out<=0;
   48788: out<=1;
   48789: out<=1;
   48790: out<=0;
   48791: out<=0;
   48792: out<=1;
   48793: out<=1;
   48794: out<=1;
   48795: out<=1;
   48796: out<=1;
   48797: out<=0;
   48798: out<=0;
   48799: out<=1;
   48800: out<=0;
   48801: out<=1;
   48802: out<=1;
   48803: out<=0;
   48804: out<=0;
   48805: out<=0;
   48806: out<=0;
   48807: out<=0;
   48808: out<=1;
   48809: out<=1;
   48810: out<=0;
   48811: out<=0;
   48812: out<=1;
   48813: out<=0;
   48814: out<=1;
   48815: out<=0;
   48816: out<=1;
   48817: out<=1;
   48818: out<=1;
   48819: out<=1;
   48820: out<=0;
   48821: out<=1;
   48822: out<=1;
   48823: out<=0;
   48824: out<=1;
   48825: out<=0;
   48826: out<=1;
   48827: out<=0;
   48828: out<=0;
   48829: out<=0;
   48830: out<=1;
   48831: out<=1;
   48832: out<=1;
   48833: out<=1;
   48834: out<=0;
   48835: out<=0;
   48836: out<=0;
   48837: out<=1;
   48838: out<=0;
   48839: out<=1;
   48840: out<=0;
   48841: out<=1;
   48842: out<=1;
   48843: out<=0;
   48844: out<=1;
   48845: out<=1;
   48846: out<=1;
   48847: out<=1;
   48848: out<=1;
   48849: out<=0;
   48850: out<=1;
   48851: out<=0;
   48852: out<=1;
   48853: out<=1;
   48854: out<=0;
   48855: out<=0;
   48856: out<=1;
   48857: out<=1;
   48858: out<=1;
   48859: out<=1;
   48860: out<=1;
   48861: out<=0;
   48862: out<=0;
   48863: out<=1;
   48864: out<=0;
   48865: out<=1;
   48866: out<=1;
   48867: out<=0;
   48868: out<=0;
   48869: out<=0;
   48870: out<=0;
   48871: out<=0;
   48872: out<=1;
   48873: out<=1;
   48874: out<=0;
   48875: out<=0;
   48876: out<=1;
   48877: out<=0;
   48878: out<=1;
   48879: out<=0;
   48880: out<=0;
   48881: out<=0;
   48882: out<=0;
   48883: out<=0;
   48884: out<=1;
   48885: out<=0;
   48886: out<=0;
   48887: out<=1;
   48888: out<=0;
   48889: out<=1;
   48890: out<=0;
   48891: out<=1;
   48892: out<=1;
   48893: out<=1;
   48894: out<=0;
   48895: out<=0;
   48896: out<=1;
   48897: out<=0;
   48898: out<=1;
   48899: out<=0;
   48900: out<=1;
   48901: out<=1;
   48902: out<=0;
   48903: out<=0;
   48904: out<=1;
   48905: out<=1;
   48906: out<=1;
   48907: out<=1;
   48908: out<=1;
   48909: out<=0;
   48910: out<=0;
   48911: out<=1;
   48912: out<=0;
   48913: out<=0;
   48914: out<=1;
   48915: out<=1;
   48916: out<=1;
   48917: out<=0;
   48918: out<=1;
   48919: out<=0;
   48920: out<=1;
   48921: out<=0;
   48922: out<=0;
   48923: out<=1;
   48924: out<=0;
   48925: out<=0;
   48926: out<=0;
   48927: out<=0;
   48928: out<=0;
   48929: out<=0;
   48930: out<=0;
   48931: out<=0;
   48932: out<=1;
   48933: out<=0;
   48934: out<=0;
   48935: out<=1;
   48936: out<=0;
   48937: out<=1;
   48938: out<=0;
   48939: out<=1;
   48940: out<=1;
   48941: out<=1;
   48942: out<=0;
   48943: out<=0;
   48944: out<=1;
   48945: out<=0;
   48946: out<=0;
   48947: out<=1;
   48948: out<=1;
   48949: out<=1;
   48950: out<=1;
   48951: out<=1;
   48952: out<=0;
   48953: out<=0;
   48954: out<=1;
   48955: out<=1;
   48956: out<=0;
   48957: out<=1;
   48958: out<=0;
   48959: out<=1;
   48960: out<=1;
   48961: out<=0;
   48962: out<=1;
   48963: out<=0;
   48964: out<=1;
   48965: out<=1;
   48966: out<=0;
   48967: out<=0;
   48968: out<=1;
   48969: out<=1;
   48970: out<=1;
   48971: out<=1;
   48972: out<=1;
   48973: out<=0;
   48974: out<=0;
   48975: out<=1;
   48976: out<=1;
   48977: out<=1;
   48978: out<=0;
   48979: out<=0;
   48980: out<=0;
   48981: out<=1;
   48982: out<=0;
   48983: out<=1;
   48984: out<=0;
   48985: out<=1;
   48986: out<=1;
   48987: out<=0;
   48988: out<=1;
   48989: out<=1;
   48990: out<=1;
   48991: out<=1;
   48992: out<=1;
   48993: out<=1;
   48994: out<=1;
   48995: out<=1;
   48996: out<=0;
   48997: out<=1;
   48998: out<=1;
   48999: out<=0;
   49000: out<=1;
   49001: out<=0;
   49002: out<=1;
   49003: out<=0;
   49004: out<=0;
   49005: out<=0;
   49006: out<=1;
   49007: out<=1;
   49008: out<=1;
   49009: out<=0;
   49010: out<=0;
   49011: out<=1;
   49012: out<=1;
   49013: out<=1;
   49014: out<=1;
   49015: out<=1;
   49016: out<=0;
   49017: out<=0;
   49018: out<=1;
   49019: out<=1;
   49020: out<=0;
   49021: out<=1;
   49022: out<=0;
   49023: out<=1;
   49024: out<=1;
   49025: out<=0;
   49026: out<=1;
   49027: out<=0;
   49028: out<=1;
   49029: out<=1;
   49030: out<=0;
   49031: out<=0;
   49032: out<=1;
   49033: out<=1;
   49034: out<=1;
   49035: out<=1;
   49036: out<=1;
   49037: out<=0;
   49038: out<=0;
   49039: out<=1;
   49040: out<=1;
   49041: out<=1;
   49042: out<=0;
   49043: out<=0;
   49044: out<=0;
   49045: out<=1;
   49046: out<=0;
   49047: out<=1;
   49048: out<=0;
   49049: out<=1;
   49050: out<=1;
   49051: out<=0;
   49052: out<=1;
   49053: out<=1;
   49054: out<=1;
   49055: out<=1;
   49056: out<=0;
   49057: out<=0;
   49058: out<=0;
   49059: out<=0;
   49060: out<=1;
   49061: out<=0;
   49062: out<=0;
   49063: out<=1;
   49064: out<=0;
   49065: out<=1;
   49066: out<=0;
   49067: out<=1;
   49068: out<=1;
   49069: out<=1;
   49070: out<=0;
   49071: out<=0;
   49072: out<=0;
   49073: out<=1;
   49074: out<=1;
   49075: out<=0;
   49076: out<=0;
   49077: out<=0;
   49078: out<=0;
   49079: out<=0;
   49080: out<=1;
   49081: out<=1;
   49082: out<=0;
   49083: out<=0;
   49084: out<=1;
   49085: out<=0;
   49086: out<=1;
   49087: out<=0;
   49088: out<=1;
   49089: out<=0;
   49090: out<=1;
   49091: out<=0;
   49092: out<=1;
   49093: out<=1;
   49094: out<=0;
   49095: out<=0;
   49096: out<=1;
   49097: out<=1;
   49098: out<=1;
   49099: out<=1;
   49100: out<=1;
   49101: out<=0;
   49102: out<=0;
   49103: out<=1;
   49104: out<=0;
   49105: out<=0;
   49106: out<=1;
   49107: out<=1;
   49108: out<=1;
   49109: out<=0;
   49110: out<=1;
   49111: out<=0;
   49112: out<=1;
   49113: out<=0;
   49114: out<=0;
   49115: out<=1;
   49116: out<=0;
   49117: out<=0;
   49118: out<=0;
   49119: out<=0;
   49120: out<=1;
   49121: out<=1;
   49122: out<=1;
   49123: out<=1;
   49124: out<=0;
   49125: out<=1;
   49126: out<=1;
   49127: out<=0;
   49128: out<=1;
   49129: out<=0;
   49130: out<=1;
   49131: out<=0;
   49132: out<=0;
   49133: out<=0;
   49134: out<=1;
   49135: out<=1;
   49136: out<=0;
   49137: out<=1;
   49138: out<=1;
   49139: out<=0;
   49140: out<=0;
   49141: out<=0;
   49142: out<=0;
   49143: out<=0;
   49144: out<=1;
   49145: out<=1;
   49146: out<=0;
   49147: out<=0;
   49148: out<=1;
   49149: out<=0;
   49150: out<=1;
   49151: out<=0;
   49152: out<=1;
   49153: out<=0;
   49154: out<=1;
   49155: out<=0;
   49156: out<=1;
   49157: out<=1;
   49158: out<=0;
   49159: out<=0;
   49160: out<=1;
   49161: out<=1;
   49162: out<=1;
   49163: out<=1;
   49164: out<=1;
   49165: out<=0;
   49166: out<=0;
   49167: out<=1;
   49168: out<=0;
   49169: out<=0;
   49170: out<=1;
   49171: out<=1;
   49172: out<=1;
   49173: out<=0;
   49174: out<=1;
   49175: out<=0;
   49176: out<=1;
   49177: out<=0;
   49178: out<=0;
   49179: out<=1;
   49180: out<=0;
   49181: out<=0;
   49182: out<=0;
   49183: out<=0;
   49184: out<=1;
   49185: out<=1;
   49186: out<=1;
   49187: out<=1;
   49188: out<=0;
   49189: out<=1;
   49190: out<=1;
   49191: out<=0;
   49192: out<=1;
   49193: out<=0;
   49194: out<=1;
   49195: out<=0;
   49196: out<=0;
   49197: out<=0;
   49198: out<=1;
   49199: out<=1;
   49200: out<=0;
   49201: out<=1;
   49202: out<=1;
   49203: out<=0;
   49204: out<=0;
   49205: out<=0;
   49206: out<=0;
   49207: out<=0;
   49208: out<=1;
   49209: out<=1;
   49210: out<=0;
   49211: out<=0;
   49212: out<=1;
   49213: out<=0;
   49214: out<=1;
   49215: out<=0;
   49216: out<=0;
   49217: out<=1;
   49218: out<=0;
   49219: out<=1;
   49220: out<=0;
   49221: out<=0;
   49222: out<=1;
   49223: out<=1;
   49224: out<=0;
   49225: out<=0;
   49226: out<=0;
   49227: out<=0;
   49228: out<=0;
   49229: out<=1;
   49230: out<=1;
   49231: out<=0;
   49232: out<=0;
   49233: out<=0;
   49234: out<=1;
   49235: out<=1;
   49236: out<=1;
   49237: out<=0;
   49238: out<=1;
   49239: out<=0;
   49240: out<=1;
   49241: out<=0;
   49242: out<=0;
   49243: out<=1;
   49244: out<=0;
   49245: out<=0;
   49246: out<=0;
   49247: out<=0;
   49248: out<=1;
   49249: out<=1;
   49250: out<=1;
   49251: out<=1;
   49252: out<=0;
   49253: out<=1;
   49254: out<=1;
   49255: out<=0;
   49256: out<=1;
   49257: out<=0;
   49258: out<=1;
   49259: out<=0;
   49260: out<=0;
   49261: out<=0;
   49262: out<=1;
   49263: out<=1;
   49264: out<=1;
   49265: out<=0;
   49266: out<=0;
   49267: out<=1;
   49268: out<=1;
   49269: out<=1;
   49270: out<=1;
   49271: out<=1;
   49272: out<=0;
   49273: out<=0;
   49274: out<=1;
   49275: out<=1;
   49276: out<=0;
   49277: out<=1;
   49278: out<=0;
   49279: out<=1;
   49280: out<=0;
   49281: out<=1;
   49282: out<=0;
   49283: out<=1;
   49284: out<=0;
   49285: out<=0;
   49286: out<=1;
   49287: out<=1;
   49288: out<=0;
   49289: out<=0;
   49290: out<=0;
   49291: out<=0;
   49292: out<=0;
   49293: out<=1;
   49294: out<=1;
   49295: out<=0;
   49296: out<=0;
   49297: out<=0;
   49298: out<=1;
   49299: out<=1;
   49300: out<=1;
   49301: out<=0;
   49302: out<=1;
   49303: out<=0;
   49304: out<=1;
   49305: out<=0;
   49306: out<=0;
   49307: out<=1;
   49308: out<=0;
   49309: out<=0;
   49310: out<=0;
   49311: out<=0;
   49312: out<=0;
   49313: out<=0;
   49314: out<=0;
   49315: out<=0;
   49316: out<=1;
   49317: out<=0;
   49318: out<=0;
   49319: out<=1;
   49320: out<=0;
   49321: out<=1;
   49322: out<=0;
   49323: out<=1;
   49324: out<=1;
   49325: out<=1;
   49326: out<=0;
   49327: out<=0;
   49328: out<=0;
   49329: out<=1;
   49330: out<=1;
   49331: out<=0;
   49332: out<=0;
   49333: out<=0;
   49334: out<=0;
   49335: out<=0;
   49336: out<=1;
   49337: out<=1;
   49338: out<=0;
   49339: out<=0;
   49340: out<=1;
   49341: out<=0;
   49342: out<=1;
   49343: out<=0;
   49344: out<=1;
   49345: out<=0;
   49346: out<=1;
   49347: out<=0;
   49348: out<=1;
   49349: out<=1;
   49350: out<=0;
   49351: out<=0;
   49352: out<=1;
   49353: out<=1;
   49354: out<=1;
   49355: out<=1;
   49356: out<=1;
   49357: out<=0;
   49358: out<=0;
   49359: out<=1;
   49360: out<=0;
   49361: out<=0;
   49362: out<=1;
   49363: out<=1;
   49364: out<=1;
   49365: out<=0;
   49366: out<=1;
   49367: out<=0;
   49368: out<=1;
   49369: out<=0;
   49370: out<=0;
   49371: out<=1;
   49372: out<=0;
   49373: out<=0;
   49374: out<=0;
   49375: out<=0;
   49376: out<=0;
   49377: out<=0;
   49378: out<=0;
   49379: out<=0;
   49380: out<=1;
   49381: out<=0;
   49382: out<=0;
   49383: out<=1;
   49384: out<=0;
   49385: out<=1;
   49386: out<=0;
   49387: out<=1;
   49388: out<=1;
   49389: out<=1;
   49390: out<=0;
   49391: out<=0;
   49392: out<=1;
   49393: out<=0;
   49394: out<=0;
   49395: out<=1;
   49396: out<=1;
   49397: out<=1;
   49398: out<=1;
   49399: out<=1;
   49400: out<=0;
   49401: out<=0;
   49402: out<=1;
   49403: out<=1;
   49404: out<=0;
   49405: out<=1;
   49406: out<=0;
   49407: out<=1;
   49408: out<=0;
   49409: out<=0;
   49410: out<=1;
   49411: out<=1;
   49412: out<=1;
   49413: out<=0;
   49414: out<=1;
   49415: out<=0;
   49416: out<=1;
   49417: out<=0;
   49418: out<=0;
   49419: out<=1;
   49420: out<=0;
   49421: out<=0;
   49422: out<=0;
   49423: out<=0;
   49424: out<=0;
   49425: out<=1;
   49426: out<=0;
   49427: out<=1;
   49428: out<=0;
   49429: out<=0;
   49430: out<=1;
   49431: out<=1;
   49432: out<=0;
   49433: out<=0;
   49434: out<=0;
   49435: out<=0;
   49436: out<=0;
   49437: out<=1;
   49438: out<=1;
   49439: out<=0;
   49440: out<=1;
   49441: out<=0;
   49442: out<=0;
   49443: out<=1;
   49444: out<=1;
   49445: out<=1;
   49446: out<=1;
   49447: out<=1;
   49448: out<=0;
   49449: out<=0;
   49450: out<=1;
   49451: out<=1;
   49452: out<=0;
   49453: out<=1;
   49454: out<=0;
   49455: out<=1;
   49456: out<=1;
   49457: out<=1;
   49458: out<=1;
   49459: out<=1;
   49460: out<=0;
   49461: out<=1;
   49462: out<=1;
   49463: out<=0;
   49464: out<=1;
   49465: out<=0;
   49466: out<=1;
   49467: out<=0;
   49468: out<=0;
   49469: out<=0;
   49470: out<=1;
   49471: out<=1;
   49472: out<=0;
   49473: out<=0;
   49474: out<=1;
   49475: out<=1;
   49476: out<=1;
   49477: out<=0;
   49478: out<=1;
   49479: out<=0;
   49480: out<=1;
   49481: out<=0;
   49482: out<=0;
   49483: out<=1;
   49484: out<=0;
   49485: out<=0;
   49486: out<=0;
   49487: out<=0;
   49488: out<=1;
   49489: out<=0;
   49490: out<=1;
   49491: out<=0;
   49492: out<=1;
   49493: out<=1;
   49494: out<=0;
   49495: out<=0;
   49496: out<=1;
   49497: out<=1;
   49498: out<=1;
   49499: out<=1;
   49500: out<=1;
   49501: out<=0;
   49502: out<=0;
   49503: out<=1;
   49504: out<=0;
   49505: out<=1;
   49506: out<=1;
   49507: out<=0;
   49508: out<=0;
   49509: out<=0;
   49510: out<=0;
   49511: out<=0;
   49512: out<=1;
   49513: out<=1;
   49514: out<=0;
   49515: out<=0;
   49516: out<=1;
   49517: out<=0;
   49518: out<=1;
   49519: out<=0;
   49520: out<=1;
   49521: out<=1;
   49522: out<=1;
   49523: out<=1;
   49524: out<=0;
   49525: out<=1;
   49526: out<=1;
   49527: out<=0;
   49528: out<=1;
   49529: out<=0;
   49530: out<=1;
   49531: out<=0;
   49532: out<=0;
   49533: out<=0;
   49534: out<=1;
   49535: out<=1;
   49536: out<=0;
   49537: out<=0;
   49538: out<=1;
   49539: out<=1;
   49540: out<=1;
   49541: out<=0;
   49542: out<=1;
   49543: out<=0;
   49544: out<=1;
   49545: out<=0;
   49546: out<=0;
   49547: out<=1;
   49548: out<=0;
   49549: out<=0;
   49550: out<=0;
   49551: out<=0;
   49552: out<=1;
   49553: out<=0;
   49554: out<=1;
   49555: out<=0;
   49556: out<=1;
   49557: out<=1;
   49558: out<=0;
   49559: out<=0;
   49560: out<=1;
   49561: out<=1;
   49562: out<=1;
   49563: out<=1;
   49564: out<=1;
   49565: out<=0;
   49566: out<=0;
   49567: out<=1;
   49568: out<=1;
   49569: out<=0;
   49570: out<=0;
   49571: out<=1;
   49572: out<=1;
   49573: out<=1;
   49574: out<=1;
   49575: out<=1;
   49576: out<=0;
   49577: out<=0;
   49578: out<=1;
   49579: out<=1;
   49580: out<=0;
   49581: out<=1;
   49582: out<=0;
   49583: out<=1;
   49584: out<=0;
   49585: out<=0;
   49586: out<=0;
   49587: out<=0;
   49588: out<=1;
   49589: out<=0;
   49590: out<=0;
   49591: out<=1;
   49592: out<=0;
   49593: out<=1;
   49594: out<=0;
   49595: out<=1;
   49596: out<=1;
   49597: out<=1;
   49598: out<=0;
   49599: out<=0;
   49600: out<=0;
   49601: out<=0;
   49602: out<=1;
   49603: out<=1;
   49604: out<=1;
   49605: out<=0;
   49606: out<=1;
   49607: out<=0;
   49608: out<=1;
   49609: out<=0;
   49610: out<=0;
   49611: out<=1;
   49612: out<=0;
   49613: out<=0;
   49614: out<=0;
   49615: out<=0;
   49616: out<=0;
   49617: out<=1;
   49618: out<=0;
   49619: out<=1;
   49620: out<=0;
   49621: out<=0;
   49622: out<=1;
   49623: out<=1;
   49624: out<=0;
   49625: out<=0;
   49626: out<=0;
   49627: out<=0;
   49628: out<=0;
   49629: out<=1;
   49630: out<=1;
   49631: out<=0;
   49632: out<=0;
   49633: out<=1;
   49634: out<=1;
   49635: out<=0;
   49636: out<=0;
   49637: out<=0;
   49638: out<=0;
   49639: out<=0;
   49640: out<=1;
   49641: out<=1;
   49642: out<=0;
   49643: out<=0;
   49644: out<=1;
   49645: out<=0;
   49646: out<=1;
   49647: out<=0;
   49648: out<=0;
   49649: out<=0;
   49650: out<=0;
   49651: out<=0;
   49652: out<=1;
   49653: out<=0;
   49654: out<=0;
   49655: out<=1;
   49656: out<=0;
   49657: out<=1;
   49658: out<=0;
   49659: out<=1;
   49660: out<=1;
   49661: out<=1;
   49662: out<=0;
   49663: out<=0;
   49664: out<=0;
   49665: out<=0;
   49666: out<=0;
   49667: out<=0;
   49668: out<=1;
   49669: out<=0;
   49670: out<=0;
   49671: out<=1;
   49672: out<=0;
   49673: out<=1;
   49674: out<=0;
   49675: out<=1;
   49676: out<=1;
   49677: out<=1;
   49678: out<=0;
   49679: out<=0;
   49680: out<=0;
   49681: out<=1;
   49682: out<=1;
   49683: out<=0;
   49684: out<=0;
   49685: out<=0;
   49686: out<=0;
   49687: out<=0;
   49688: out<=1;
   49689: out<=1;
   49690: out<=0;
   49691: out<=0;
   49692: out<=1;
   49693: out<=0;
   49694: out<=1;
   49695: out<=0;
   49696: out<=0;
   49697: out<=1;
   49698: out<=0;
   49699: out<=1;
   49700: out<=0;
   49701: out<=0;
   49702: out<=1;
   49703: out<=1;
   49704: out<=0;
   49705: out<=0;
   49706: out<=0;
   49707: out<=0;
   49708: out<=0;
   49709: out<=1;
   49710: out<=1;
   49711: out<=0;
   49712: out<=0;
   49713: out<=0;
   49714: out<=1;
   49715: out<=1;
   49716: out<=1;
   49717: out<=0;
   49718: out<=1;
   49719: out<=0;
   49720: out<=1;
   49721: out<=0;
   49722: out<=0;
   49723: out<=1;
   49724: out<=0;
   49725: out<=0;
   49726: out<=0;
   49727: out<=0;
   49728: out<=0;
   49729: out<=0;
   49730: out<=0;
   49731: out<=0;
   49732: out<=1;
   49733: out<=0;
   49734: out<=0;
   49735: out<=1;
   49736: out<=0;
   49737: out<=1;
   49738: out<=0;
   49739: out<=1;
   49740: out<=1;
   49741: out<=1;
   49742: out<=0;
   49743: out<=0;
   49744: out<=1;
   49745: out<=0;
   49746: out<=0;
   49747: out<=1;
   49748: out<=1;
   49749: out<=1;
   49750: out<=1;
   49751: out<=1;
   49752: out<=0;
   49753: out<=0;
   49754: out<=1;
   49755: out<=1;
   49756: out<=0;
   49757: out<=1;
   49758: out<=0;
   49759: out<=1;
   49760: out<=1;
   49761: out<=0;
   49762: out<=1;
   49763: out<=0;
   49764: out<=1;
   49765: out<=1;
   49766: out<=0;
   49767: out<=0;
   49768: out<=1;
   49769: out<=1;
   49770: out<=1;
   49771: out<=1;
   49772: out<=1;
   49773: out<=0;
   49774: out<=0;
   49775: out<=1;
   49776: out<=0;
   49777: out<=0;
   49778: out<=1;
   49779: out<=1;
   49780: out<=1;
   49781: out<=0;
   49782: out<=1;
   49783: out<=0;
   49784: out<=1;
   49785: out<=0;
   49786: out<=0;
   49787: out<=1;
   49788: out<=0;
   49789: out<=0;
   49790: out<=0;
   49791: out<=0;
   49792: out<=1;
   49793: out<=1;
   49794: out<=1;
   49795: out<=1;
   49796: out<=0;
   49797: out<=1;
   49798: out<=1;
   49799: out<=0;
   49800: out<=1;
   49801: out<=0;
   49802: out<=1;
   49803: out<=0;
   49804: out<=0;
   49805: out<=0;
   49806: out<=1;
   49807: out<=1;
   49808: out<=0;
   49809: out<=1;
   49810: out<=1;
   49811: out<=0;
   49812: out<=0;
   49813: out<=0;
   49814: out<=0;
   49815: out<=0;
   49816: out<=1;
   49817: out<=1;
   49818: out<=0;
   49819: out<=0;
   49820: out<=1;
   49821: out<=0;
   49822: out<=1;
   49823: out<=0;
   49824: out<=1;
   49825: out<=0;
   49826: out<=1;
   49827: out<=0;
   49828: out<=1;
   49829: out<=1;
   49830: out<=0;
   49831: out<=0;
   49832: out<=1;
   49833: out<=1;
   49834: out<=1;
   49835: out<=1;
   49836: out<=1;
   49837: out<=0;
   49838: out<=0;
   49839: out<=1;
   49840: out<=0;
   49841: out<=0;
   49842: out<=1;
   49843: out<=1;
   49844: out<=1;
   49845: out<=0;
   49846: out<=1;
   49847: out<=0;
   49848: out<=1;
   49849: out<=0;
   49850: out<=0;
   49851: out<=1;
   49852: out<=0;
   49853: out<=0;
   49854: out<=0;
   49855: out<=0;
   49856: out<=1;
   49857: out<=1;
   49858: out<=1;
   49859: out<=1;
   49860: out<=0;
   49861: out<=1;
   49862: out<=1;
   49863: out<=0;
   49864: out<=1;
   49865: out<=0;
   49866: out<=1;
   49867: out<=0;
   49868: out<=0;
   49869: out<=0;
   49870: out<=1;
   49871: out<=1;
   49872: out<=1;
   49873: out<=0;
   49874: out<=0;
   49875: out<=1;
   49876: out<=1;
   49877: out<=1;
   49878: out<=1;
   49879: out<=1;
   49880: out<=0;
   49881: out<=0;
   49882: out<=1;
   49883: out<=1;
   49884: out<=0;
   49885: out<=1;
   49886: out<=0;
   49887: out<=1;
   49888: out<=0;
   49889: out<=1;
   49890: out<=0;
   49891: out<=1;
   49892: out<=0;
   49893: out<=0;
   49894: out<=1;
   49895: out<=1;
   49896: out<=0;
   49897: out<=0;
   49898: out<=0;
   49899: out<=0;
   49900: out<=0;
   49901: out<=1;
   49902: out<=1;
   49903: out<=0;
   49904: out<=0;
   49905: out<=0;
   49906: out<=1;
   49907: out<=1;
   49908: out<=1;
   49909: out<=0;
   49910: out<=1;
   49911: out<=0;
   49912: out<=1;
   49913: out<=0;
   49914: out<=0;
   49915: out<=1;
   49916: out<=0;
   49917: out<=0;
   49918: out<=0;
   49919: out<=0;
   49920: out<=1;
   49921: out<=0;
   49922: out<=0;
   49923: out<=1;
   49924: out<=1;
   49925: out<=1;
   49926: out<=1;
   49927: out<=1;
   49928: out<=0;
   49929: out<=0;
   49930: out<=1;
   49931: out<=1;
   49932: out<=0;
   49933: out<=1;
   49934: out<=0;
   49935: out<=1;
   49936: out<=0;
   49937: out<=0;
   49938: out<=0;
   49939: out<=0;
   49940: out<=1;
   49941: out<=0;
   49942: out<=0;
   49943: out<=1;
   49944: out<=0;
   49945: out<=1;
   49946: out<=0;
   49947: out<=1;
   49948: out<=1;
   49949: out<=1;
   49950: out<=0;
   49951: out<=0;
   49952: out<=0;
   49953: out<=0;
   49954: out<=1;
   49955: out<=1;
   49956: out<=1;
   49957: out<=0;
   49958: out<=1;
   49959: out<=0;
   49960: out<=1;
   49961: out<=0;
   49962: out<=0;
   49963: out<=1;
   49964: out<=0;
   49965: out<=0;
   49966: out<=0;
   49967: out<=0;
   49968: out<=1;
   49969: out<=0;
   49970: out<=1;
   49971: out<=0;
   49972: out<=1;
   49973: out<=1;
   49974: out<=0;
   49975: out<=0;
   49976: out<=1;
   49977: out<=1;
   49978: out<=1;
   49979: out<=1;
   49980: out<=1;
   49981: out<=0;
   49982: out<=0;
   49983: out<=1;
   49984: out<=0;
   49985: out<=1;
   49986: out<=1;
   49987: out<=0;
   49988: out<=0;
   49989: out<=0;
   49990: out<=0;
   49991: out<=0;
   49992: out<=1;
   49993: out<=1;
   49994: out<=0;
   49995: out<=0;
   49996: out<=1;
   49997: out<=0;
   49998: out<=1;
   49999: out<=0;
   50000: out<=0;
   50001: out<=0;
   50002: out<=0;
   50003: out<=0;
   50004: out<=1;
   50005: out<=0;
   50006: out<=0;
   50007: out<=1;
   50008: out<=0;
   50009: out<=1;
   50010: out<=0;
   50011: out<=1;
   50012: out<=1;
   50013: out<=1;
   50014: out<=0;
   50015: out<=0;
   50016: out<=0;
   50017: out<=0;
   50018: out<=1;
   50019: out<=1;
   50020: out<=1;
   50021: out<=0;
   50022: out<=1;
   50023: out<=0;
   50024: out<=1;
   50025: out<=0;
   50026: out<=0;
   50027: out<=1;
   50028: out<=0;
   50029: out<=0;
   50030: out<=0;
   50031: out<=0;
   50032: out<=0;
   50033: out<=1;
   50034: out<=0;
   50035: out<=1;
   50036: out<=0;
   50037: out<=0;
   50038: out<=1;
   50039: out<=1;
   50040: out<=0;
   50041: out<=0;
   50042: out<=0;
   50043: out<=0;
   50044: out<=0;
   50045: out<=1;
   50046: out<=1;
   50047: out<=0;
   50048: out<=1;
   50049: out<=0;
   50050: out<=0;
   50051: out<=1;
   50052: out<=1;
   50053: out<=1;
   50054: out<=1;
   50055: out<=1;
   50056: out<=0;
   50057: out<=0;
   50058: out<=1;
   50059: out<=1;
   50060: out<=0;
   50061: out<=1;
   50062: out<=0;
   50063: out<=1;
   50064: out<=1;
   50065: out<=1;
   50066: out<=1;
   50067: out<=1;
   50068: out<=0;
   50069: out<=1;
   50070: out<=1;
   50071: out<=0;
   50072: out<=1;
   50073: out<=0;
   50074: out<=1;
   50075: out<=0;
   50076: out<=0;
   50077: out<=0;
   50078: out<=1;
   50079: out<=1;
   50080: out<=0;
   50081: out<=0;
   50082: out<=1;
   50083: out<=1;
   50084: out<=1;
   50085: out<=0;
   50086: out<=1;
   50087: out<=0;
   50088: out<=1;
   50089: out<=0;
   50090: out<=0;
   50091: out<=1;
   50092: out<=0;
   50093: out<=0;
   50094: out<=0;
   50095: out<=0;
   50096: out<=0;
   50097: out<=1;
   50098: out<=0;
   50099: out<=1;
   50100: out<=0;
   50101: out<=0;
   50102: out<=1;
   50103: out<=1;
   50104: out<=0;
   50105: out<=0;
   50106: out<=0;
   50107: out<=0;
   50108: out<=0;
   50109: out<=1;
   50110: out<=1;
   50111: out<=0;
   50112: out<=0;
   50113: out<=1;
   50114: out<=1;
   50115: out<=0;
   50116: out<=0;
   50117: out<=0;
   50118: out<=0;
   50119: out<=0;
   50120: out<=1;
   50121: out<=1;
   50122: out<=0;
   50123: out<=0;
   50124: out<=1;
   50125: out<=0;
   50126: out<=1;
   50127: out<=0;
   50128: out<=1;
   50129: out<=1;
   50130: out<=1;
   50131: out<=1;
   50132: out<=0;
   50133: out<=1;
   50134: out<=1;
   50135: out<=0;
   50136: out<=1;
   50137: out<=0;
   50138: out<=1;
   50139: out<=0;
   50140: out<=0;
   50141: out<=0;
   50142: out<=1;
   50143: out<=1;
   50144: out<=0;
   50145: out<=0;
   50146: out<=1;
   50147: out<=1;
   50148: out<=1;
   50149: out<=0;
   50150: out<=1;
   50151: out<=0;
   50152: out<=1;
   50153: out<=0;
   50154: out<=0;
   50155: out<=1;
   50156: out<=0;
   50157: out<=0;
   50158: out<=0;
   50159: out<=0;
   50160: out<=1;
   50161: out<=0;
   50162: out<=1;
   50163: out<=0;
   50164: out<=1;
   50165: out<=1;
   50166: out<=0;
   50167: out<=0;
   50168: out<=1;
   50169: out<=1;
   50170: out<=1;
   50171: out<=1;
   50172: out<=1;
   50173: out<=0;
   50174: out<=0;
   50175: out<=1;
   50176: out<=0;
   50177: out<=0;
   50178: out<=1;
   50179: out<=1;
   50180: out<=0;
   50181: out<=1;
   50182: out<=0;
   50183: out<=1;
   50184: out<=0;
   50185: out<=1;
   50186: out<=1;
   50187: out<=0;
   50188: out<=0;
   50189: out<=0;
   50190: out<=0;
   50191: out<=0;
   50192: out<=1;
   50193: out<=0;
   50194: out<=1;
   50195: out<=0;
   50196: out<=0;
   50197: out<=0;
   50198: out<=1;
   50199: out<=1;
   50200: out<=0;
   50201: out<=0;
   50202: out<=0;
   50203: out<=0;
   50204: out<=1;
   50205: out<=0;
   50206: out<=0;
   50207: out<=1;
   50208: out<=0;
   50209: out<=1;
   50210: out<=1;
   50211: out<=0;
   50212: out<=1;
   50213: out<=1;
   50214: out<=1;
   50215: out<=1;
   50216: out<=0;
   50217: out<=0;
   50218: out<=1;
   50219: out<=1;
   50220: out<=1;
   50221: out<=0;
   50222: out<=1;
   50223: out<=0;
   50224: out<=1;
   50225: out<=1;
   50226: out<=1;
   50227: out<=1;
   50228: out<=1;
   50229: out<=0;
   50230: out<=0;
   50231: out<=1;
   50232: out<=0;
   50233: out<=1;
   50234: out<=0;
   50235: out<=1;
   50236: out<=0;
   50237: out<=0;
   50238: out<=1;
   50239: out<=1;
   50240: out<=0;
   50241: out<=0;
   50242: out<=1;
   50243: out<=1;
   50244: out<=0;
   50245: out<=1;
   50246: out<=0;
   50247: out<=1;
   50248: out<=0;
   50249: out<=1;
   50250: out<=1;
   50251: out<=0;
   50252: out<=0;
   50253: out<=0;
   50254: out<=0;
   50255: out<=0;
   50256: out<=0;
   50257: out<=1;
   50258: out<=0;
   50259: out<=1;
   50260: out<=1;
   50261: out<=1;
   50262: out<=0;
   50263: out<=0;
   50264: out<=1;
   50265: out<=1;
   50266: out<=1;
   50267: out<=1;
   50268: out<=0;
   50269: out<=1;
   50270: out<=1;
   50271: out<=0;
   50272: out<=1;
   50273: out<=0;
   50274: out<=0;
   50275: out<=1;
   50276: out<=0;
   50277: out<=0;
   50278: out<=0;
   50279: out<=0;
   50280: out<=1;
   50281: out<=1;
   50282: out<=0;
   50283: out<=0;
   50284: out<=0;
   50285: out<=1;
   50286: out<=0;
   50287: out<=1;
   50288: out<=1;
   50289: out<=1;
   50290: out<=1;
   50291: out<=1;
   50292: out<=1;
   50293: out<=0;
   50294: out<=0;
   50295: out<=1;
   50296: out<=0;
   50297: out<=1;
   50298: out<=0;
   50299: out<=1;
   50300: out<=0;
   50301: out<=0;
   50302: out<=1;
   50303: out<=1;
   50304: out<=0;
   50305: out<=0;
   50306: out<=1;
   50307: out<=1;
   50308: out<=0;
   50309: out<=1;
   50310: out<=0;
   50311: out<=1;
   50312: out<=0;
   50313: out<=1;
   50314: out<=1;
   50315: out<=0;
   50316: out<=0;
   50317: out<=0;
   50318: out<=0;
   50319: out<=0;
   50320: out<=0;
   50321: out<=1;
   50322: out<=0;
   50323: out<=1;
   50324: out<=1;
   50325: out<=1;
   50326: out<=0;
   50327: out<=0;
   50328: out<=1;
   50329: out<=1;
   50330: out<=1;
   50331: out<=1;
   50332: out<=0;
   50333: out<=1;
   50334: out<=1;
   50335: out<=0;
   50336: out<=0;
   50337: out<=1;
   50338: out<=1;
   50339: out<=0;
   50340: out<=1;
   50341: out<=1;
   50342: out<=1;
   50343: out<=1;
   50344: out<=0;
   50345: out<=0;
   50346: out<=1;
   50347: out<=1;
   50348: out<=1;
   50349: out<=0;
   50350: out<=1;
   50351: out<=0;
   50352: out<=0;
   50353: out<=0;
   50354: out<=0;
   50355: out<=0;
   50356: out<=0;
   50357: out<=1;
   50358: out<=1;
   50359: out<=0;
   50360: out<=1;
   50361: out<=0;
   50362: out<=1;
   50363: out<=0;
   50364: out<=1;
   50365: out<=1;
   50366: out<=0;
   50367: out<=0;
   50368: out<=0;
   50369: out<=0;
   50370: out<=1;
   50371: out<=1;
   50372: out<=0;
   50373: out<=1;
   50374: out<=0;
   50375: out<=1;
   50376: out<=0;
   50377: out<=1;
   50378: out<=1;
   50379: out<=0;
   50380: out<=0;
   50381: out<=0;
   50382: out<=0;
   50383: out<=0;
   50384: out<=1;
   50385: out<=0;
   50386: out<=1;
   50387: out<=0;
   50388: out<=0;
   50389: out<=0;
   50390: out<=1;
   50391: out<=1;
   50392: out<=0;
   50393: out<=0;
   50394: out<=0;
   50395: out<=0;
   50396: out<=1;
   50397: out<=0;
   50398: out<=0;
   50399: out<=1;
   50400: out<=1;
   50401: out<=0;
   50402: out<=0;
   50403: out<=1;
   50404: out<=0;
   50405: out<=0;
   50406: out<=0;
   50407: out<=0;
   50408: out<=1;
   50409: out<=1;
   50410: out<=0;
   50411: out<=0;
   50412: out<=0;
   50413: out<=1;
   50414: out<=0;
   50415: out<=1;
   50416: out<=0;
   50417: out<=0;
   50418: out<=0;
   50419: out<=0;
   50420: out<=0;
   50421: out<=1;
   50422: out<=1;
   50423: out<=0;
   50424: out<=1;
   50425: out<=0;
   50426: out<=1;
   50427: out<=0;
   50428: out<=1;
   50429: out<=1;
   50430: out<=0;
   50431: out<=0;
   50432: out<=0;
   50433: out<=1;
   50434: out<=0;
   50435: out<=1;
   50436: out<=1;
   50437: out<=1;
   50438: out<=0;
   50439: out<=0;
   50440: out<=1;
   50441: out<=1;
   50442: out<=1;
   50443: out<=1;
   50444: out<=0;
   50445: out<=1;
   50446: out<=1;
   50447: out<=0;
   50448: out<=0;
   50449: out<=0;
   50450: out<=1;
   50451: out<=1;
   50452: out<=0;
   50453: out<=1;
   50454: out<=0;
   50455: out<=1;
   50456: out<=0;
   50457: out<=1;
   50458: out<=1;
   50459: out<=0;
   50460: out<=0;
   50461: out<=0;
   50462: out<=0;
   50463: out<=0;
   50464: out<=1;
   50465: out<=1;
   50466: out<=1;
   50467: out<=1;
   50468: out<=1;
   50469: out<=0;
   50470: out<=0;
   50471: out<=1;
   50472: out<=0;
   50473: out<=1;
   50474: out<=0;
   50475: out<=1;
   50476: out<=0;
   50477: out<=0;
   50478: out<=1;
   50479: out<=1;
   50480: out<=1;
   50481: out<=0;
   50482: out<=0;
   50483: out<=1;
   50484: out<=0;
   50485: out<=0;
   50486: out<=0;
   50487: out<=0;
   50488: out<=1;
   50489: out<=1;
   50490: out<=0;
   50491: out<=0;
   50492: out<=0;
   50493: out<=1;
   50494: out<=0;
   50495: out<=1;
   50496: out<=1;
   50497: out<=0;
   50498: out<=1;
   50499: out<=0;
   50500: out<=0;
   50501: out<=0;
   50502: out<=1;
   50503: out<=1;
   50504: out<=0;
   50505: out<=0;
   50506: out<=0;
   50507: out<=0;
   50508: out<=1;
   50509: out<=0;
   50510: out<=0;
   50511: out<=1;
   50512: out<=0;
   50513: out<=0;
   50514: out<=1;
   50515: out<=1;
   50516: out<=0;
   50517: out<=1;
   50518: out<=0;
   50519: out<=1;
   50520: out<=0;
   50521: out<=1;
   50522: out<=1;
   50523: out<=0;
   50524: out<=0;
   50525: out<=0;
   50526: out<=0;
   50527: out<=0;
   50528: out<=1;
   50529: out<=1;
   50530: out<=1;
   50531: out<=1;
   50532: out<=1;
   50533: out<=0;
   50534: out<=0;
   50535: out<=1;
   50536: out<=0;
   50537: out<=1;
   50538: out<=0;
   50539: out<=1;
   50540: out<=0;
   50541: out<=0;
   50542: out<=1;
   50543: out<=1;
   50544: out<=0;
   50545: out<=1;
   50546: out<=1;
   50547: out<=0;
   50548: out<=1;
   50549: out<=1;
   50550: out<=1;
   50551: out<=1;
   50552: out<=0;
   50553: out<=0;
   50554: out<=1;
   50555: out<=1;
   50556: out<=1;
   50557: out<=0;
   50558: out<=1;
   50559: out<=0;
   50560: out<=1;
   50561: out<=0;
   50562: out<=1;
   50563: out<=0;
   50564: out<=0;
   50565: out<=0;
   50566: out<=1;
   50567: out<=1;
   50568: out<=0;
   50569: out<=0;
   50570: out<=0;
   50571: out<=0;
   50572: out<=1;
   50573: out<=0;
   50574: out<=0;
   50575: out<=1;
   50576: out<=0;
   50577: out<=0;
   50578: out<=1;
   50579: out<=1;
   50580: out<=0;
   50581: out<=1;
   50582: out<=0;
   50583: out<=1;
   50584: out<=0;
   50585: out<=1;
   50586: out<=1;
   50587: out<=0;
   50588: out<=0;
   50589: out<=0;
   50590: out<=0;
   50591: out<=0;
   50592: out<=0;
   50593: out<=0;
   50594: out<=0;
   50595: out<=0;
   50596: out<=0;
   50597: out<=1;
   50598: out<=1;
   50599: out<=0;
   50600: out<=1;
   50601: out<=0;
   50602: out<=1;
   50603: out<=0;
   50604: out<=1;
   50605: out<=1;
   50606: out<=0;
   50607: out<=0;
   50608: out<=1;
   50609: out<=0;
   50610: out<=0;
   50611: out<=1;
   50612: out<=0;
   50613: out<=0;
   50614: out<=0;
   50615: out<=0;
   50616: out<=1;
   50617: out<=1;
   50618: out<=0;
   50619: out<=0;
   50620: out<=0;
   50621: out<=1;
   50622: out<=0;
   50623: out<=1;
   50624: out<=0;
   50625: out<=1;
   50626: out<=0;
   50627: out<=1;
   50628: out<=1;
   50629: out<=1;
   50630: out<=0;
   50631: out<=0;
   50632: out<=1;
   50633: out<=1;
   50634: out<=1;
   50635: out<=1;
   50636: out<=0;
   50637: out<=1;
   50638: out<=1;
   50639: out<=0;
   50640: out<=0;
   50641: out<=0;
   50642: out<=1;
   50643: out<=1;
   50644: out<=0;
   50645: out<=1;
   50646: out<=0;
   50647: out<=1;
   50648: out<=0;
   50649: out<=1;
   50650: out<=1;
   50651: out<=0;
   50652: out<=0;
   50653: out<=0;
   50654: out<=0;
   50655: out<=0;
   50656: out<=0;
   50657: out<=0;
   50658: out<=0;
   50659: out<=0;
   50660: out<=0;
   50661: out<=1;
   50662: out<=1;
   50663: out<=0;
   50664: out<=1;
   50665: out<=0;
   50666: out<=1;
   50667: out<=0;
   50668: out<=1;
   50669: out<=1;
   50670: out<=0;
   50671: out<=0;
   50672: out<=0;
   50673: out<=1;
   50674: out<=1;
   50675: out<=0;
   50676: out<=1;
   50677: out<=1;
   50678: out<=1;
   50679: out<=1;
   50680: out<=0;
   50681: out<=0;
   50682: out<=1;
   50683: out<=1;
   50684: out<=1;
   50685: out<=0;
   50686: out<=1;
   50687: out<=0;
   50688: out<=0;
   50689: out<=1;
   50690: out<=1;
   50691: out<=0;
   50692: out<=1;
   50693: out<=1;
   50694: out<=1;
   50695: out<=1;
   50696: out<=0;
   50697: out<=0;
   50698: out<=1;
   50699: out<=1;
   50700: out<=1;
   50701: out<=0;
   50702: out<=1;
   50703: out<=0;
   50704: out<=0;
   50705: out<=0;
   50706: out<=0;
   50707: out<=0;
   50708: out<=0;
   50709: out<=1;
   50710: out<=1;
   50711: out<=0;
   50712: out<=1;
   50713: out<=0;
   50714: out<=1;
   50715: out<=0;
   50716: out<=1;
   50717: out<=1;
   50718: out<=0;
   50719: out<=0;
   50720: out<=0;
   50721: out<=0;
   50722: out<=1;
   50723: out<=1;
   50724: out<=0;
   50725: out<=1;
   50726: out<=0;
   50727: out<=1;
   50728: out<=0;
   50729: out<=1;
   50730: out<=1;
   50731: out<=0;
   50732: out<=0;
   50733: out<=0;
   50734: out<=0;
   50735: out<=0;
   50736: out<=0;
   50737: out<=1;
   50738: out<=0;
   50739: out<=1;
   50740: out<=1;
   50741: out<=1;
   50742: out<=0;
   50743: out<=0;
   50744: out<=1;
   50745: out<=1;
   50746: out<=1;
   50747: out<=1;
   50748: out<=0;
   50749: out<=1;
   50750: out<=1;
   50751: out<=0;
   50752: out<=1;
   50753: out<=0;
   50754: out<=0;
   50755: out<=1;
   50756: out<=0;
   50757: out<=0;
   50758: out<=0;
   50759: out<=0;
   50760: out<=1;
   50761: out<=1;
   50762: out<=0;
   50763: out<=0;
   50764: out<=0;
   50765: out<=1;
   50766: out<=0;
   50767: out<=1;
   50768: out<=0;
   50769: out<=0;
   50770: out<=0;
   50771: out<=0;
   50772: out<=0;
   50773: out<=1;
   50774: out<=1;
   50775: out<=0;
   50776: out<=1;
   50777: out<=0;
   50778: out<=1;
   50779: out<=0;
   50780: out<=1;
   50781: out<=1;
   50782: out<=0;
   50783: out<=0;
   50784: out<=0;
   50785: out<=0;
   50786: out<=1;
   50787: out<=1;
   50788: out<=0;
   50789: out<=1;
   50790: out<=0;
   50791: out<=1;
   50792: out<=0;
   50793: out<=1;
   50794: out<=1;
   50795: out<=0;
   50796: out<=0;
   50797: out<=0;
   50798: out<=0;
   50799: out<=0;
   50800: out<=1;
   50801: out<=0;
   50802: out<=1;
   50803: out<=0;
   50804: out<=0;
   50805: out<=0;
   50806: out<=1;
   50807: out<=1;
   50808: out<=0;
   50809: out<=0;
   50810: out<=0;
   50811: out<=0;
   50812: out<=1;
   50813: out<=0;
   50814: out<=0;
   50815: out<=1;
   50816: out<=0;
   50817: out<=1;
   50818: out<=1;
   50819: out<=0;
   50820: out<=1;
   50821: out<=1;
   50822: out<=1;
   50823: out<=1;
   50824: out<=0;
   50825: out<=0;
   50826: out<=1;
   50827: out<=1;
   50828: out<=1;
   50829: out<=0;
   50830: out<=1;
   50831: out<=0;
   50832: out<=1;
   50833: out<=1;
   50834: out<=1;
   50835: out<=1;
   50836: out<=1;
   50837: out<=0;
   50838: out<=0;
   50839: out<=1;
   50840: out<=0;
   50841: out<=1;
   50842: out<=0;
   50843: out<=1;
   50844: out<=0;
   50845: out<=0;
   50846: out<=1;
   50847: out<=1;
   50848: out<=0;
   50849: out<=0;
   50850: out<=1;
   50851: out<=1;
   50852: out<=0;
   50853: out<=1;
   50854: out<=0;
   50855: out<=1;
   50856: out<=0;
   50857: out<=1;
   50858: out<=1;
   50859: out<=0;
   50860: out<=0;
   50861: out<=0;
   50862: out<=0;
   50863: out<=0;
   50864: out<=1;
   50865: out<=0;
   50866: out<=1;
   50867: out<=0;
   50868: out<=0;
   50869: out<=0;
   50870: out<=1;
   50871: out<=1;
   50872: out<=0;
   50873: out<=0;
   50874: out<=0;
   50875: out<=0;
   50876: out<=1;
   50877: out<=0;
   50878: out<=0;
   50879: out<=1;
   50880: out<=1;
   50881: out<=0;
   50882: out<=0;
   50883: out<=1;
   50884: out<=0;
   50885: out<=0;
   50886: out<=0;
   50887: out<=0;
   50888: out<=1;
   50889: out<=1;
   50890: out<=0;
   50891: out<=0;
   50892: out<=0;
   50893: out<=1;
   50894: out<=0;
   50895: out<=1;
   50896: out<=1;
   50897: out<=1;
   50898: out<=1;
   50899: out<=1;
   50900: out<=1;
   50901: out<=0;
   50902: out<=0;
   50903: out<=1;
   50904: out<=0;
   50905: out<=1;
   50906: out<=0;
   50907: out<=1;
   50908: out<=0;
   50909: out<=0;
   50910: out<=1;
   50911: out<=1;
   50912: out<=0;
   50913: out<=0;
   50914: out<=1;
   50915: out<=1;
   50916: out<=0;
   50917: out<=1;
   50918: out<=0;
   50919: out<=1;
   50920: out<=0;
   50921: out<=1;
   50922: out<=1;
   50923: out<=0;
   50924: out<=0;
   50925: out<=0;
   50926: out<=0;
   50927: out<=0;
   50928: out<=0;
   50929: out<=1;
   50930: out<=0;
   50931: out<=1;
   50932: out<=1;
   50933: out<=1;
   50934: out<=0;
   50935: out<=0;
   50936: out<=1;
   50937: out<=1;
   50938: out<=1;
   50939: out<=1;
   50940: out<=0;
   50941: out<=1;
   50942: out<=1;
   50943: out<=0;
   50944: out<=0;
   50945: out<=0;
   50946: out<=0;
   50947: out<=0;
   50948: out<=0;
   50949: out<=1;
   50950: out<=1;
   50951: out<=0;
   50952: out<=1;
   50953: out<=0;
   50954: out<=1;
   50955: out<=0;
   50956: out<=1;
   50957: out<=1;
   50958: out<=0;
   50959: out<=0;
   50960: out<=1;
   50961: out<=0;
   50962: out<=0;
   50963: out<=1;
   50964: out<=0;
   50965: out<=0;
   50966: out<=0;
   50967: out<=0;
   50968: out<=1;
   50969: out<=1;
   50970: out<=0;
   50971: out<=0;
   50972: out<=0;
   50973: out<=1;
   50974: out<=0;
   50975: out<=1;
   50976: out<=1;
   50977: out<=0;
   50978: out<=1;
   50979: out<=0;
   50980: out<=0;
   50981: out<=0;
   50982: out<=1;
   50983: out<=1;
   50984: out<=0;
   50985: out<=0;
   50986: out<=0;
   50987: out<=0;
   50988: out<=1;
   50989: out<=0;
   50990: out<=0;
   50991: out<=1;
   50992: out<=0;
   50993: out<=0;
   50994: out<=1;
   50995: out<=1;
   50996: out<=0;
   50997: out<=1;
   50998: out<=0;
   50999: out<=1;
   51000: out<=0;
   51001: out<=1;
   51002: out<=1;
   51003: out<=0;
   51004: out<=0;
   51005: out<=0;
   51006: out<=0;
   51007: out<=0;
   51008: out<=0;
   51009: out<=0;
   51010: out<=0;
   51011: out<=0;
   51012: out<=0;
   51013: out<=1;
   51014: out<=1;
   51015: out<=0;
   51016: out<=1;
   51017: out<=0;
   51018: out<=1;
   51019: out<=0;
   51020: out<=1;
   51021: out<=1;
   51022: out<=0;
   51023: out<=0;
   51024: out<=0;
   51025: out<=1;
   51026: out<=1;
   51027: out<=0;
   51028: out<=1;
   51029: out<=1;
   51030: out<=1;
   51031: out<=1;
   51032: out<=0;
   51033: out<=0;
   51034: out<=1;
   51035: out<=1;
   51036: out<=1;
   51037: out<=0;
   51038: out<=1;
   51039: out<=0;
   51040: out<=0;
   51041: out<=1;
   51042: out<=0;
   51043: out<=1;
   51044: out<=1;
   51045: out<=1;
   51046: out<=0;
   51047: out<=0;
   51048: out<=1;
   51049: out<=1;
   51050: out<=1;
   51051: out<=1;
   51052: out<=0;
   51053: out<=1;
   51054: out<=1;
   51055: out<=0;
   51056: out<=0;
   51057: out<=0;
   51058: out<=1;
   51059: out<=1;
   51060: out<=0;
   51061: out<=1;
   51062: out<=0;
   51063: out<=1;
   51064: out<=0;
   51065: out<=1;
   51066: out<=1;
   51067: out<=0;
   51068: out<=0;
   51069: out<=0;
   51070: out<=0;
   51071: out<=0;
   51072: out<=1;
   51073: out<=1;
   51074: out<=1;
   51075: out<=1;
   51076: out<=1;
   51077: out<=0;
   51078: out<=0;
   51079: out<=1;
   51080: out<=0;
   51081: out<=1;
   51082: out<=0;
   51083: out<=1;
   51084: out<=0;
   51085: out<=0;
   51086: out<=1;
   51087: out<=1;
   51088: out<=1;
   51089: out<=0;
   51090: out<=0;
   51091: out<=1;
   51092: out<=0;
   51093: out<=0;
   51094: out<=0;
   51095: out<=0;
   51096: out<=1;
   51097: out<=1;
   51098: out<=0;
   51099: out<=0;
   51100: out<=0;
   51101: out<=1;
   51102: out<=0;
   51103: out<=1;
   51104: out<=0;
   51105: out<=1;
   51106: out<=0;
   51107: out<=1;
   51108: out<=1;
   51109: out<=1;
   51110: out<=0;
   51111: out<=0;
   51112: out<=1;
   51113: out<=1;
   51114: out<=1;
   51115: out<=1;
   51116: out<=0;
   51117: out<=1;
   51118: out<=1;
   51119: out<=0;
   51120: out<=0;
   51121: out<=0;
   51122: out<=1;
   51123: out<=1;
   51124: out<=0;
   51125: out<=1;
   51126: out<=0;
   51127: out<=1;
   51128: out<=0;
   51129: out<=1;
   51130: out<=1;
   51131: out<=0;
   51132: out<=0;
   51133: out<=0;
   51134: out<=0;
   51135: out<=0;
   51136: out<=1;
   51137: out<=1;
   51138: out<=1;
   51139: out<=1;
   51140: out<=1;
   51141: out<=0;
   51142: out<=0;
   51143: out<=1;
   51144: out<=0;
   51145: out<=1;
   51146: out<=0;
   51147: out<=1;
   51148: out<=0;
   51149: out<=0;
   51150: out<=1;
   51151: out<=1;
   51152: out<=0;
   51153: out<=1;
   51154: out<=1;
   51155: out<=0;
   51156: out<=1;
   51157: out<=1;
   51158: out<=1;
   51159: out<=1;
   51160: out<=0;
   51161: out<=0;
   51162: out<=1;
   51163: out<=1;
   51164: out<=1;
   51165: out<=0;
   51166: out<=1;
   51167: out<=0;
   51168: out<=1;
   51169: out<=0;
   51170: out<=1;
   51171: out<=0;
   51172: out<=0;
   51173: out<=0;
   51174: out<=1;
   51175: out<=1;
   51176: out<=0;
   51177: out<=0;
   51178: out<=0;
   51179: out<=0;
   51180: out<=1;
   51181: out<=0;
   51182: out<=0;
   51183: out<=1;
   51184: out<=0;
   51185: out<=0;
   51186: out<=1;
   51187: out<=1;
   51188: out<=0;
   51189: out<=1;
   51190: out<=0;
   51191: out<=1;
   51192: out<=0;
   51193: out<=1;
   51194: out<=1;
   51195: out<=0;
   51196: out<=0;
   51197: out<=0;
   51198: out<=0;
   51199: out<=0;
   51200: out<=0;
   51201: out<=0;
   51202: out<=0;
   51203: out<=0;
   51204: out<=0;
   51205: out<=1;
   51206: out<=1;
   51207: out<=0;
   51208: out<=0;
   51209: out<=1;
   51210: out<=0;
   51211: out<=1;
   51212: out<=0;
   51213: out<=0;
   51214: out<=1;
   51215: out<=1;
   51216: out<=1;
   51217: out<=0;
   51218: out<=0;
   51219: out<=1;
   51220: out<=0;
   51221: out<=0;
   51222: out<=0;
   51223: out<=0;
   51224: out<=0;
   51225: out<=0;
   51226: out<=1;
   51227: out<=1;
   51228: out<=1;
   51229: out<=0;
   51230: out<=1;
   51231: out<=0;
   51232: out<=0;
   51233: out<=1;
   51234: out<=0;
   51235: out<=1;
   51236: out<=1;
   51237: out<=1;
   51238: out<=0;
   51239: out<=0;
   51240: out<=0;
   51241: out<=0;
   51242: out<=0;
   51243: out<=0;
   51244: out<=1;
   51245: out<=0;
   51246: out<=0;
   51247: out<=1;
   51248: out<=1;
   51249: out<=1;
   51250: out<=0;
   51251: out<=0;
   51252: out<=1;
   51253: out<=0;
   51254: out<=1;
   51255: out<=0;
   51256: out<=0;
   51257: out<=1;
   51258: out<=1;
   51259: out<=0;
   51260: out<=0;
   51261: out<=0;
   51262: out<=0;
   51263: out<=0;
   51264: out<=0;
   51265: out<=0;
   51266: out<=0;
   51267: out<=0;
   51268: out<=0;
   51269: out<=1;
   51270: out<=1;
   51271: out<=0;
   51272: out<=0;
   51273: out<=1;
   51274: out<=0;
   51275: out<=1;
   51276: out<=0;
   51277: out<=0;
   51278: out<=1;
   51279: out<=1;
   51280: out<=0;
   51281: out<=1;
   51282: out<=1;
   51283: out<=0;
   51284: out<=1;
   51285: out<=1;
   51286: out<=1;
   51287: out<=1;
   51288: out<=1;
   51289: out<=1;
   51290: out<=0;
   51291: out<=0;
   51292: out<=0;
   51293: out<=1;
   51294: out<=0;
   51295: out<=1;
   51296: out<=1;
   51297: out<=0;
   51298: out<=1;
   51299: out<=0;
   51300: out<=0;
   51301: out<=0;
   51302: out<=1;
   51303: out<=1;
   51304: out<=1;
   51305: out<=1;
   51306: out<=1;
   51307: out<=1;
   51308: out<=0;
   51309: out<=1;
   51310: out<=1;
   51311: out<=0;
   51312: out<=1;
   51313: out<=1;
   51314: out<=0;
   51315: out<=0;
   51316: out<=1;
   51317: out<=0;
   51318: out<=1;
   51319: out<=0;
   51320: out<=0;
   51321: out<=1;
   51322: out<=1;
   51323: out<=0;
   51324: out<=0;
   51325: out<=0;
   51326: out<=0;
   51327: out<=0;
   51328: out<=1;
   51329: out<=1;
   51330: out<=1;
   51331: out<=1;
   51332: out<=1;
   51333: out<=0;
   51334: out<=0;
   51335: out<=1;
   51336: out<=1;
   51337: out<=0;
   51338: out<=1;
   51339: out<=0;
   51340: out<=1;
   51341: out<=1;
   51342: out<=0;
   51343: out<=0;
   51344: out<=1;
   51345: out<=0;
   51346: out<=0;
   51347: out<=1;
   51348: out<=0;
   51349: out<=0;
   51350: out<=0;
   51351: out<=0;
   51352: out<=0;
   51353: out<=0;
   51354: out<=1;
   51355: out<=1;
   51356: out<=1;
   51357: out<=0;
   51358: out<=1;
   51359: out<=0;
   51360: out<=1;
   51361: out<=0;
   51362: out<=1;
   51363: out<=0;
   51364: out<=0;
   51365: out<=0;
   51366: out<=1;
   51367: out<=1;
   51368: out<=1;
   51369: out<=1;
   51370: out<=1;
   51371: out<=1;
   51372: out<=0;
   51373: out<=1;
   51374: out<=1;
   51375: out<=0;
   51376: out<=1;
   51377: out<=1;
   51378: out<=0;
   51379: out<=0;
   51380: out<=1;
   51381: out<=0;
   51382: out<=1;
   51383: out<=0;
   51384: out<=0;
   51385: out<=1;
   51386: out<=1;
   51387: out<=0;
   51388: out<=0;
   51389: out<=0;
   51390: out<=0;
   51391: out<=0;
   51392: out<=1;
   51393: out<=1;
   51394: out<=1;
   51395: out<=1;
   51396: out<=1;
   51397: out<=0;
   51398: out<=0;
   51399: out<=1;
   51400: out<=1;
   51401: out<=0;
   51402: out<=1;
   51403: out<=0;
   51404: out<=1;
   51405: out<=1;
   51406: out<=0;
   51407: out<=0;
   51408: out<=0;
   51409: out<=1;
   51410: out<=1;
   51411: out<=0;
   51412: out<=1;
   51413: out<=1;
   51414: out<=1;
   51415: out<=1;
   51416: out<=1;
   51417: out<=1;
   51418: out<=0;
   51419: out<=0;
   51420: out<=0;
   51421: out<=1;
   51422: out<=0;
   51423: out<=1;
   51424: out<=0;
   51425: out<=1;
   51426: out<=0;
   51427: out<=1;
   51428: out<=1;
   51429: out<=1;
   51430: out<=0;
   51431: out<=0;
   51432: out<=0;
   51433: out<=0;
   51434: out<=0;
   51435: out<=0;
   51436: out<=1;
   51437: out<=0;
   51438: out<=0;
   51439: out<=1;
   51440: out<=1;
   51441: out<=1;
   51442: out<=0;
   51443: out<=0;
   51444: out<=1;
   51445: out<=0;
   51446: out<=1;
   51447: out<=0;
   51448: out<=0;
   51449: out<=1;
   51450: out<=1;
   51451: out<=0;
   51452: out<=0;
   51453: out<=0;
   51454: out<=0;
   51455: out<=0;
   51456: out<=0;
   51457: out<=1;
   51458: out<=1;
   51459: out<=0;
   51460: out<=1;
   51461: out<=1;
   51462: out<=1;
   51463: out<=1;
   51464: out<=1;
   51465: out<=1;
   51466: out<=0;
   51467: out<=0;
   51468: out<=0;
   51469: out<=1;
   51470: out<=0;
   51471: out<=1;
   51472: out<=0;
   51473: out<=0;
   51474: out<=0;
   51475: out<=0;
   51476: out<=0;
   51477: out<=1;
   51478: out<=1;
   51479: out<=0;
   51480: out<=0;
   51481: out<=1;
   51482: out<=0;
   51483: out<=1;
   51484: out<=0;
   51485: out<=0;
   51486: out<=1;
   51487: out<=1;
   51488: out<=1;
   51489: out<=1;
   51490: out<=0;
   51491: out<=0;
   51492: out<=1;
   51493: out<=0;
   51494: out<=1;
   51495: out<=0;
   51496: out<=0;
   51497: out<=1;
   51498: out<=1;
   51499: out<=0;
   51500: out<=0;
   51501: out<=0;
   51502: out<=0;
   51503: out<=0;
   51504: out<=1;
   51505: out<=0;
   51506: out<=1;
   51507: out<=0;
   51508: out<=0;
   51509: out<=0;
   51510: out<=1;
   51511: out<=1;
   51512: out<=1;
   51513: out<=1;
   51514: out<=1;
   51515: out<=1;
   51516: out<=0;
   51517: out<=1;
   51518: out<=1;
   51519: out<=0;
   51520: out<=1;
   51521: out<=0;
   51522: out<=0;
   51523: out<=1;
   51524: out<=0;
   51525: out<=0;
   51526: out<=0;
   51527: out<=0;
   51528: out<=0;
   51529: out<=0;
   51530: out<=1;
   51531: out<=1;
   51532: out<=1;
   51533: out<=0;
   51534: out<=1;
   51535: out<=0;
   51536: out<=0;
   51537: out<=0;
   51538: out<=0;
   51539: out<=0;
   51540: out<=0;
   51541: out<=1;
   51542: out<=1;
   51543: out<=0;
   51544: out<=0;
   51545: out<=1;
   51546: out<=0;
   51547: out<=1;
   51548: out<=0;
   51549: out<=0;
   51550: out<=1;
   51551: out<=1;
   51552: out<=1;
   51553: out<=1;
   51554: out<=0;
   51555: out<=0;
   51556: out<=1;
   51557: out<=0;
   51558: out<=1;
   51559: out<=0;
   51560: out<=0;
   51561: out<=1;
   51562: out<=1;
   51563: out<=0;
   51564: out<=0;
   51565: out<=0;
   51566: out<=0;
   51567: out<=0;
   51568: out<=0;
   51569: out<=1;
   51570: out<=0;
   51571: out<=1;
   51572: out<=1;
   51573: out<=1;
   51574: out<=0;
   51575: out<=0;
   51576: out<=0;
   51577: out<=0;
   51578: out<=0;
   51579: out<=0;
   51580: out<=1;
   51581: out<=0;
   51582: out<=0;
   51583: out<=1;
   51584: out<=0;
   51585: out<=1;
   51586: out<=1;
   51587: out<=0;
   51588: out<=1;
   51589: out<=1;
   51590: out<=1;
   51591: out<=1;
   51592: out<=1;
   51593: out<=1;
   51594: out<=0;
   51595: out<=0;
   51596: out<=0;
   51597: out<=1;
   51598: out<=0;
   51599: out<=1;
   51600: out<=1;
   51601: out<=1;
   51602: out<=1;
   51603: out<=1;
   51604: out<=1;
   51605: out<=0;
   51606: out<=0;
   51607: out<=1;
   51608: out<=1;
   51609: out<=0;
   51610: out<=1;
   51611: out<=0;
   51612: out<=1;
   51613: out<=1;
   51614: out<=0;
   51615: out<=0;
   51616: out<=1;
   51617: out<=1;
   51618: out<=0;
   51619: out<=0;
   51620: out<=1;
   51621: out<=0;
   51622: out<=1;
   51623: out<=0;
   51624: out<=0;
   51625: out<=1;
   51626: out<=1;
   51627: out<=0;
   51628: out<=0;
   51629: out<=0;
   51630: out<=0;
   51631: out<=0;
   51632: out<=0;
   51633: out<=1;
   51634: out<=0;
   51635: out<=1;
   51636: out<=1;
   51637: out<=1;
   51638: out<=0;
   51639: out<=0;
   51640: out<=0;
   51641: out<=0;
   51642: out<=0;
   51643: out<=0;
   51644: out<=1;
   51645: out<=0;
   51646: out<=0;
   51647: out<=1;
   51648: out<=1;
   51649: out<=0;
   51650: out<=0;
   51651: out<=1;
   51652: out<=0;
   51653: out<=0;
   51654: out<=0;
   51655: out<=0;
   51656: out<=0;
   51657: out<=0;
   51658: out<=1;
   51659: out<=1;
   51660: out<=1;
   51661: out<=0;
   51662: out<=1;
   51663: out<=0;
   51664: out<=1;
   51665: out<=1;
   51666: out<=1;
   51667: out<=1;
   51668: out<=1;
   51669: out<=0;
   51670: out<=0;
   51671: out<=1;
   51672: out<=1;
   51673: out<=0;
   51674: out<=1;
   51675: out<=0;
   51676: out<=1;
   51677: out<=1;
   51678: out<=0;
   51679: out<=0;
   51680: out<=1;
   51681: out<=1;
   51682: out<=0;
   51683: out<=0;
   51684: out<=1;
   51685: out<=0;
   51686: out<=1;
   51687: out<=0;
   51688: out<=0;
   51689: out<=1;
   51690: out<=1;
   51691: out<=0;
   51692: out<=0;
   51693: out<=0;
   51694: out<=0;
   51695: out<=0;
   51696: out<=1;
   51697: out<=0;
   51698: out<=1;
   51699: out<=0;
   51700: out<=0;
   51701: out<=0;
   51702: out<=1;
   51703: out<=1;
   51704: out<=1;
   51705: out<=1;
   51706: out<=1;
   51707: out<=1;
   51708: out<=0;
   51709: out<=1;
   51710: out<=1;
   51711: out<=0;
   51712: out<=1;
   51713: out<=0;
   51714: out<=1;
   51715: out<=0;
   51716: out<=0;
   51717: out<=0;
   51718: out<=1;
   51719: out<=1;
   51720: out<=1;
   51721: out<=1;
   51722: out<=1;
   51723: out<=1;
   51724: out<=0;
   51725: out<=1;
   51726: out<=1;
   51727: out<=0;
   51728: out<=1;
   51729: out<=1;
   51730: out<=0;
   51731: out<=0;
   51732: out<=1;
   51733: out<=0;
   51734: out<=1;
   51735: out<=0;
   51736: out<=0;
   51737: out<=1;
   51738: out<=1;
   51739: out<=0;
   51740: out<=0;
   51741: out<=0;
   51742: out<=0;
   51743: out<=0;
   51744: out<=1;
   51745: out<=1;
   51746: out<=1;
   51747: out<=1;
   51748: out<=1;
   51749: out<=0;
   51750: out<=0;
   51751: out<=1;
   51752: out<=1;
   51753: out<=0;
   51754: out<=1;
   51755: out<=0;
   51756: out<=1;
   51757: out<=1;
   51758: out<=0;
   51759: out<=0;
   51760: out<=1;
   51761: out<=0;
   51762: out<=0;
   51763: out<=1;
   51764: out<=0;
   51765: out<=0;
   51766: out<=0;
   51767: out<=0;
   51768: out<=0;
   51769: out<=0;
   51770: out<=1;
   51771: out<=1;
   51772: out<=1;
   51773: out<=0;
   51774: out<=1;
   51775: out<=0;
   51776: out<=0;
   51777: out<=1;
   51778: out<=0;
   51779: out<=1;
   51780: out<=1;
   51781: out<=1;
   51782: out<=0;
   51783: out<=0;
   51784: out<=0;
   51785: out<=0;
   51786: out<=0;
   51787: out<=0;
   51788: out<=1;
   51789: out<=0;
   51790: out<=0;
   51791: out<=1;
   51792: out<=1;
   51793: out<=1;
   51794: out<=0;
   51795: out<=0;
   51796: out<=1;
   51797: out<=0;
   51798: out<=1;
   51799: out<=0;
   51800: out<=0;
   51801: out<=1;
   51802: out<=1;
   51803: out<=0;
   51804: out<=0;
   51805: out<=0;
   51806: out<=0;
   51807: out<=0;
   51808: out<=1;
   51809: out<=1;
   51810: out<=1;
   51811: out<=1;
   51812: out<=1;
   51813: out<=0;
   51814: out<=0;
   51815: out<=1;
   51816: out<=1;
   51817: out<=0;
   51818: out<=1;
   51819: out<=0;
   51820: out<=1;
   51821: out<=1;
   51822: out<=0;
   51823: out<=0;
   51824: out<=0;
   51825: out<=1;
   51826: out<=1;
   51827: out<=0;
   51828: out<=1;
   51829: out<=1;
   51830: out<=1;
   51831: out<=1;
   51832: out<=1;
   51833: out<=1;
   51834: out<=0;
   51835: out<=0;
   51836: out<=0;
   51837: out<=1;
   51838: out<=0;
   51839: out<=1;
   51840: out<=0;
   51841: out<=1;
   51842: out<=0;
   51843: out<=1;
   51844: out<=1;
   51845: out<=1;
   51846: out<=0;
   51847: out<=0;
   51848: out<=0;
   51849: out<=0;
   51850: out<=0;
   51851: out<=0;
   51852: out<=1;
   51853: out<=0;
   51854: out<=0;
   51855: out<=1;
   51856: out<=1;
   51857: out<=1;
   51858: out<=0;
   51859: out<=0;
   51860: out<=1;
   51861: out<=0;
   51862: out<=1;
   51863: out<=0;
   51864: out<=0;
   51865: out<=1;
   51866: out<=1;
   51867: out<=0;
   51868: out<=0;
   51869: out<=0;
   51870: out<=0;
   51871: out<=0;
   51872: out<=0;
   51873: out<=0;
   51874: out<=0;
   51875: out<=0;
   51876: out<=0;
   51877: out<=1;
   51878: out<=1;
   51879: out<=0;
   51880: out<=0;
   51881: out<=1;
   51882: out<=0;
   51883: out<=1;
   51884: out<=0;
   51885: out<=0;
   51886: out<=1;
   51887: out<=1;
   51888: out<=1;
   51889: out<=0;
   51890: out<=0;
   51891: out<=1;
   51892: out<=0;
   51893: out<=0;
   51894: out<=0;
   51895: out<=0;
   51896: out<=0;
   51897: out<=0;
   51898: out<=1;
   51899: out<=1;
   51900: out<=1;
   51901: out<=0;
   51902: out<=1;
   51903: out<=0;
   51904: out<=1;
   51905: out<=0;
   51906: out<=1;
   51907: out<=0;
   51908: out<=0;
   51909: out<=0;
   51910: out<=1;
   51911: out<=1;
   51912: out<=1;
   51913: out<=1;
   51914: out<=1;
   51915: out<=1;
   51916: out<=0;
   51917: out<=1;
   51918: out<=1;
   51919: out<=0;
   51920: out<=1;
   51921: out<=1;
   51922: out<=0;
   51923: out<=0;
   51924: out<=1;
   51925: out<=0;
   51926: out<=1;
   51927: out<=0;
   51928: out<=0;
   51929: out<=1;
   51930: out<=1;
   51931: out<=0;
   51932: out<=0;
   51933: out<=0;
   51934: out<=0;
   51935: out<=0;
   51936: out<=0;
   51937: out<=0;
   51938: out<=0;
   51939: out<=0;
   51940: out<=0;
   51941: out<=1;
   51942: out<=1;
   51943: out<=0;
   51944: out<=0;
   51945: out<=1;
   51946: out<=0;
   51947: out<=1;
   51948: out<=0;
   51949: out<=0;
   51950: out<=1;
   51951: out<=1;
   51952: out<=0;
   51953: out<=1;
   51954: out<=1;
   51955: out<=0;
   51956: out<=1;
   51957: out<=1;
   51958: out<=1;
   51959: out<=1;
   51960: out<=1;
   51961: out<=1;
   51962: out<=0;
   51963: out<=0;
   51964: out<=0;
   51965: out<=1;
   51966: out<=0;
   51967: out<=1;
   51968: out<=1;
   51969: out<=1;
   51970: out<=0;
   51971: out<=0;
   51972: out<=1;
   51973: out<=0;
   51974: out<=1;
   51975: out<=0;
   51976: out<=0;
   51977: out<=1;
   51978: out<=1;
   51979: out<=0;
   51980: out<=0;
   51981: out<=0;
   51982: out<=0;
   51983: out<=0;
   51984: out<=0;
   51985: out<=1;
   51986: out<=0;
   51987: out<=1;
   51988: out<=1;
   51989: out<=1;
   51990: out<=0;
   51991: out<=0;
   51992: out<=0;
   51993: out<=0;
   51994: out<=0;
   51995: out<=0;
   51996: out<=1;
   51997: out<=0;
   51998: out<=0;
   51999: out<=1;
   52000: out<=0;
   52001: out<=1;
   52002: out<=1;
   52003: out<=0;
   52004: out<=1;
   52005: out<=1;
   52006: out<=1;
   52007: out<=1;
   52008: out<=1;
   52009: out<=1;
   52010: out<=0;
   52011: out<=0;
   52012: out<=0;
   52013: out<=1;
   52014: out<=0;
   52015: out<=1;
   52016: out<=1;
   52017: out<=1;
   52018: out<=1;
   52019: out<=1;
   52020: out<=1;
   52021: out<=0;
   52022: out<=0;
   52023: out<=1;
   52024: out<=1;
   52025: out<=0;
   52026: out<=1;
   52027: out<=0;
   52028: out<=1;
   52029: out<=1;
   52030: out<=0;
   52031: out<=0;
   52032: out<=1;
   52033: out<=1;
   52034: out<=0;
   52035: out<=0;
   52036: out<=1;
   52037: out<=0;
   52038: out<=1;
   52039: out<=0;
   52040: out<=0;
   52041: out<=1;
   52042: out<=1;
   52043: out<=0;
   52044: out<=0;
   52045: out<=0;
   52046: out<=0;
   52047: out<=0;
   52048: out<=1;
   52049: out<=0;
   52050: out<=1;
   52051: out<=0;
   52052: out<=0;
   52053: out<=0;
   52054: out<=1;
   52055: out<=1;
   52056: out<=1;
   52057: out<=1;
   52058: out<=1;
   52059: out<=1;
   52060: out<=0;
   52061: out<=1;
   52062: out<=1;
   52063: out<=0;
   52064: out<=1;
   52065: out<=0;
   52066: out<=0;
   52067: out<=1;
   52068: out<=0;
   52069: out<=0;
   52070: out<=0;
   52071: out<=0;
   52072: out<=0;
   52073: out<=0;
   52074: out<=1;
   52075: out<=1;
   52076: out<=1;
   52077: out<=0;
   52078: out<=1;
   52079: out<=0;
   52080: out<=1;
   52081: out<=1;
   52082: out<=1;
   52083: out<=1;
   52084: out<=1;
   52085: out<=0;
   52086: out<=0;
   52087: out<=1;
   52088: out<=1;
   52089: out<=0;
   52090: out<=1;
   52091: out<=0;
   52092: out<=1;
   52093: out<=1;
   52094: out<=0;
   52095: out<=0;
   52096: out<=1;
   52097: out<=1;
   52098: out<=0;
   52099: out<=0;
   52100: out<=1;
   52101: out<=0;
   52102: out<=1;
   52103: out<=0;
   52104: out<=0;
   52105: out<=1;
   52106: out<=1;
   52107: out<=0;
   52108: out<=0;
   52109: out<=0;
   52110: out<=0;
   52111: out<=0;
   52112: out<=1;
   52113: out<=0;
   52114: out<=1;
   52115: out<=0;
   52116: out<=0;
   52117: out<=0;
   52118: out<=1;
   52119: out<=1;
   52120: out<=1;
   52121: out<=1;
   52122: out<=1;
   52123: out<=1;
   52124: out<=0;
   52125: out<=1;
   52126: out<=1;
   52127: out<=0;
   52128: out<=0;
   52129: out<=1;
   52130: out<=1;
   52131: out<=0;
   52132: out<=1;
   52133: out<=1;
   52134: out<=1;
   52135: out<=1;
   52136: out<=1;
   52137: out<=1;
   52138: out<=0;
   52139: out<=0;
   52140: out<=0;
   52141: out<=1;
   52142: out<=0;
   52143: out<=1;
   52144: out<=0;
   52145: out<=0;
   52146: out<=0;
   52147: out<=0;
   52148: out<=0;
   52149: out<=1;
   52150: out<=1;
   52151: out<=0;
   52152: out<=0;
   52153: out<=1;
   52154: out<=0;
   52155: out<=1;
   52156: out<=0;
   52157: out<=0;
   52158: out<=1;
   52159: out<=1;
   52160: out<=1;
   52161: out<=1;
   52162: out<=0;
   52163: out<=0;
   52164: out<=1;
   52165: out<=0;
   52166: out<=1;
   52167: out<=0;
   52168: out<=0;
   52169: out<=1;
   52170: out<=1;
   52171: out<=0;
   52172: out<=0;
   52173: out<=0;
   52174: out<=0;
   52175: out<=0;
   52176: out<=0;
   52177: out<=1;
   52178: out<=0;
   52179: out<=1;
   52180: out<=1;
   52181: out<=1;
   52182: out<=0;
   52183: out<=0;
   52184: out<=0;
   52185: out<=0;
   52186: out<=0;
   52187: out<=0;
   52188: out<=1;
   52189: out<=0;
   52190: out<=0;
   52191: out<=1;
   52192: out<=1;
   52193: out<=0;
   52194: out<=0;
   52195: out<=1;
   52196: out<=0;
   52197: out<=0;
   52198: out<=0;
   52199: out<=0;
   52200: out<=0;
   52201: out<=0;
   52202: out<=1;
   52203: out<=1;
   52204: out<=1;
   52205: out<=0;
   52206: out<=1;
   52207: out<=0;
   52208: out<=0;
   52209: out<=0;
   52210: out<=0;
   52211: out<=0;
   52212: out<=0;
   52213: out<=1;
   52214: out<=1;
   52215: out<=0;
   52216: out<=0;
   52217: out<=1;
   52218: out<=0;
   52219: out<=1;
   52220: out<=0;
   52221: out<=0;
   52222: out<=1;
   52223: out<=1;
   52224: out<=1;
   52225: out<=0;
   52226: out<=0;
   52227: out<=1;
   52228: out<=1;
   52229: out<=1;
   52230: out<=1;
   52231: out<=1;
   52232: out<=1;
   52233: out<=1;
   52234: out<=0;
   52235: out<=0;
   52236: out<=1;
   52237: out<=0;
   52238: out<=1;
   52239: out<=0;
   52240: out<=0;
   52241: out<=0;
   52242: out<=0;
   52243: out<=0;
   52244: out<=1;
   52245: out<=0;
   52246: out<=0;
   52247: out<=1;
   52248: out<=1;
   52249: out<=0;
   52250: out<=1;
   52251: out<=0;
   52252: out<=0;
   52253: out<=0;
   52254: out<=1;
   52255: out<=1;
   52256: out<=1;
   52257: out<=1;
   52258: out<=0;
   52259: out<=0;
   52260: out<=0;
   52261: out<=1;
   52262: out<=0;
   52263: out<=1;
   52264: out<=1;
   52265: out<=0;
   52266: out<=0;
   52267: out<=1;
   52268: out<=0;
   52269: out<=0;
   52270: out<=0;
   52271: out<=0;
   52272: out<=0;
   52273: out<=1;
   52274: out<=0;
   52275: out<=1;
   52276: out<=0;
   52277: out<=0;
   52278: out<=1;
   52279: out<=1;
   52280: out<=1;
   52281: out<=1;
   52282: out<=1;
   52283: out<=1;
   52284: out<=1;
   52285: out<=0;
   52286: out<=0;
   52287: out<=1;
   52288: out<=0;
   52289: out<=1;
   52290: out<=1;
   52291: out<=0;
   52292: out<=0;
   52293: out<=0;
   52294: out<=0;
   52295: out<=0;
   52296: out<=0;
   52297: out<=0;
   52298: out<=1;
   52299: out<=1;
   52300: out<=0;
   52301: out<=1;
   52302: out<=0;
   52303: out<=1;
   52304: out<=0;
   52305: out<=0;
   52306: out<=0;
   52307: out<=0;
   52308: out<=1;
   52309: out<=0;
   52310: out<=0;
   52311: out<=1;
   52312: out<=1;
   52313: out<=0;
   52314: out<=1;
   52315: out<=0;
   52316: out<=0;
   52317: out<=0;
   52318: out<=1;
   52319: out<=1;
   52320: out<=1;
   52321: out<=1;
   52322: out<=0;
   52323: out<=0;
   52324: out<=0;
   52325: out<=1;
   52326: out<=0;
   52327: out<=1;
   52328: out<=1;
   52329: out<=0;
   52330: out<=0;
   52331: out<=1;
   52332: out<=0;
   52333: out<=0;
   52334: out<=0;
   52335: out<=0;
   52336: out<=1;
   52337: out<=0;
   52338: out<=1;
   52339: out<=0;
   52340: out<=1;
   52341: out<=1;
   52342: out<=0;
   52343: out<=0;
   52344: out<=0;
   52345: out<=0;
   52346: out<=0;
   52347: out<=0;
   52348: out<=0;
   52349: out<=1;
   52350: out<=1;
   52351: out<=0;
   52352: out<=1;
   52353: out<=0;
   52354: out<=0;
   52355: out<=1;
   52356: out<=1;
   52357: out<=1;
   52358: out<=1;
   52359: out<=1;
   52360: out<=1;
   52361: out<=1;
   52362: out<=0;
   52363: out<=0;
   52364: out<=1;
   52365: out<=0;
   52366: out<=1;
   52367: out<=0;
   52368: out<=1;
   52369: out<=1;
   52370: out<=1;
   52371: out<=1;
   52372: out<=0;
   52373: out<=1;
   52374: out<=1;
   52375: out<=0;
   52376: out<=0;
   52377: out<=1;
   52378: out<=0;
   52379: out<=1;
   52380: out<=1;
   52381: out<=1;
   52382: out<=0;
   52383: out<=0;
   52384: out<=1;
   52385: out<=1;
   52386: out<=0;
   52387: out<=0;
   52388: out<=0;
   52389: out<=1;
   52390: out<=0;
   52391: out<=1;
   52392: out<=1;
   52393: out<=0;
   52394: out<=0;
   52395: out<=1;
   52396: out<=0;
   52397: out<=0;
   52398: out<=0;
   52399: out<=0;
   52400: out<=1;
   52401: out<=0;
   52402: out<=1;
   52403: out<=0;
   52404: out<=1;
   52405: out<=1;
   52406: out<=0;
   52407: out<=0;
   52408: out<=0;
   52409: out<=0;
   52410: out<=0;
   52411: out<=0;
   52412: out<=0;
   52413: out<=1;
   52414: out<=1;
   52415: out<=0;
   52416: out<=0;
   52417: out<=1;
   52418: out<=1;
   52419: out<=0;
   52420: out<=0;
   52421: out<=0;
   52422: out<=0;
   52423: out<=0;
   52424: out<=0;
   52425: out<=0;
   52426: out<=1;
   52427: out<=1;
   52428: out<=0;
   52429: out<=1;
   52430: out<=0;
   52431: out<=1;
   52432: out<=1;
   52433: out<=1;
   52434: out<=1;
   52435: out<=1;
   52436: out<=0;
   52437: out<=1;
   52438: out<=1;
   52439: out<=0;
   52440: out<=0;
   52441: out<=1;
   52442: out<=0;
   52443: out<=1;
   52444: out<=1;
   52445: out<=1;
   52446: out<=0;
   52447: out<=0;
   52448: out<=1;
   52449: out<=1;
   52450: out<=0;
   52451: out<=0;
   52452: out<=0;
   52453: out<=1;
   52454: out<=0;
   52455: out<=1;
   52456: out<=1;
   52457: out<=0;
   52458: out<=0;
   52459: out<=1;
   52460: out<=0;
   52461: out<=0;
   52462: out<=0;
   52463: out<=0;
   52464: out<=0;
   52465: out<=1;
   52466: out<=0;
   52467: out<=1;
   52468: out<=0;
   52469: out<=0;
   52470: out<=1;
   52471: out<=1;
   52472: out<=1;
   52473: out<=1;
   52474: out<=1;
   52475: out<=1;
   52476: out<=1;
   52477: out<=0;
   52478: out<=0;
   52479: out<=1;
   52480: out<=0;
   52481: out<=0;
   52482: out<=0;
   52483: out<=0;
   52484: out<=1;
   52485: out<=0;
   52486: out<=0;
   52487: out<=1;
   52488: out<=1;
   52489: out<=0;
   52490: out<=1;
   52491: out<=0;
   52492: out<=0;
   52493: out<=0;
   52494: out<=1;
   52495: out<=1;
   52496: out<=0;
   52497: out<=1;
   52498: out<=1;
   52499: out<=0;
   52500: out<=0;
   52501: out<=0;
   52502: out<=0;
   52503: out<=0;
   52504: out<=0;
   52505: out<=0;
   52506: out<=1;
   52507: out<=1;
   52508: out<=0;
   52509: out<=1;
   52510: out<=0;
   52511: out<=1;
   52512: out<=1;
   52513: out<=0;
   52514: out<=1;
   52515: out<=0;
   52516: out<=1;
   52517: out<=1;
   52518: out<=0;
   52519: out<=0;
   52520: out<=0;
   52521: out<=0;
   52522: out<=0;
   52523: out<=0;
   52524: out<=0;
   52525: out<=1;
   52526: out<=1;
   52527: out<=0;
   52528: out<=1;
   52529: out<=1;
   52530: out<=0;
   52531: out<=0;
   52532: out<=0;
   52533: out<=1;
   52534: out<=0;
   52535: out<=1;
   52536: out<=1;
   52537: out<=0;
   52538: out<=0;
   52539: out<=1;
   52540: out<=0;
   52541: out<=0;
   52542: out<=0;
   52543: out<=0;
   52544: out<=0;
   52545: out<=0;
   52546: out<=0;
   52547: out<=0;
   52548: out<=1;
   52549: out<=0;
   52550: out<=0;
   52551: out<=1;
   52552: out<=1;
   52553: out<=0;
   52554: out<=1;
   52555: out<=0;
   52556: out<=0;
   52557: out<=0;
   52558: out<=1;
   52559: out<=1;
   52560: out<=1;
   52561: out<=0;
   52562: out<=0;
   52563: out<=1;
   52564: out<=1;
   52565: out<=1;
   52566: out<=1;
   52567: out<=1;
   52568: out<=1;
   52569: out<=1;
   52570: out<=0;
   52571: out<=0;
   52572: out<=1;
   52573: out<=0;
   52574: out<=1;
   52575: out<=0;
   52576: out<=0;
   52577: out<=1;
   52578: out<=0;
   52579: out<=1;
   52580: out<=0;
   52581: out<=0;
   52582: out<=1;
   52583: out<=1;
   52584: out<=1;
   52585: out<=1;
   52586: out<=1;
   52587: out<=1;
   52588: out<=1;
   52589: out<=0;
   52590: out<=0;
   52591: out<=1;
   52592: out<=1;
   52593: out<=1;
   52594: out<=0;
   52595: out<=0;
   52596: out<=0;
   52597: out<=1;
   52598: out<=0;
   52599: out<=1;
   52600: out<=1;
   52601: out<=0;
   52602: out<=0;
   52603: out<=1;
   52604: out<=0;
   52605: out<=0;
   52606: out<=0;
   52607: out<=0;
   52608: out<=1;
   52609: out<=1;
   52610: out<=1;
   52611: out<=1;
   52612: out<=0;
   52613: out<=1;
   52614: out<=1;
   52615: out<=0;
   52616: out<=0;
   52617: out<=1;
   52618: out<=0;
   52619: out<=1;
   52620: out<=1;
   52621: out<=1;
   52622: out<=0;
   52623: out<=0;
   52624: out<=0;
   52625: out<=1;
   52626: out<=1;
   52627: out<=0;
   52628: out<=0;
   52629: out<=0;
   52630: out<=0;
   52631: out<=0;
   52632: out<=0;
   52633: out<=0;
   52634: out<=1;
   52635: out<=1;
   52636: out<=0;
   52637: out<=1;
   52638: out<=0;
   52639: out<=1;
   52640: out<=0;
   52641: out<=1;
   52642: out<=0;
   52643: out<=1;
   52644: out<=0;
   52645: out<=0;
   52646: out<=1;
   52647: out<=1;
   52648: out<=1;
   52649: out<=1;
   52650: out<=1;
   52651: out<=1;
   52652: out<=1;
   52653: out<=0;
   52654: out<=0;
   52655: out<=1;
   52656: out<=1;
   52657: out<=1;
   52658: out<=0;
   52659: out<=0;
   52660: out<=0;
   52661: out<=1;
   52662: out<=0;
   52663: out<=1;
   52664: out<=1;
   52665: out<=0;
   52666: out<=0;
   52667: out<=1;
   52668: out<=0;
   52669: out<=0;
   52670: out<=0;
   52671: out<=0;
   52672: out<=1;
   52673: out<=1;
   52674: out<=1;
   52675: out<=1;
   52676: out<=0;
   52677: out<=1;
   52678: out<=1;
   52679: out<=0;
   52680: out<=0;
   52681: out<=1;
   52682: out<=0;
   52683: out<=1;
   52684: out<=1;
   52685: out<=1;
   52686: out<=0;
   52687: out<=0;
   52688: out<=1;
   52689: out<=0;
   52690: out<=0;
   52691: out<=1;
   52692: out<=1;
   52693: out<=1;
   52694: out<=1;
   52695: out<=1;
   52696: out<=1;
   52697: out<=1;
   52698: out<=0;
   52699: out<=0;
   52700: out<=1;
   52701: out<=0;
   52702: out<=1;
   52703: out<=0;
   52704: out<=1;
   52705: out<=0;
   52706: out<=1;
   52707: out<=0;
   52708: out<=1;
   52709: out<=1;
   52710: out<=0;
   52711: out<=0;
   52712: out<=0;
   52713: out<=0;
   52714: out<=0;
   52715: out<=0;
   52716: out<=0;
   52717: out<=1;
   52718: out<=1;
   52719: out<=0;
   52720: out<=1;
   52721: out<=1;
   52722: out<=0;
   52723: out<=0;
   52724: out<=0;
   52725: out<=1;
   52726: out<=0;
   52727: out<=1;
   52728: out<=1;
   52729: out<=0;
   52730: out<=0;
   52731: out<=1;
   52732: out<=0;
   52733: out<=0;
   52734: out<=0;
   52735: out<=0;
   52736: out<=1;
   52737: out<=1;
   52738: out<=0;
   52739: out<=0;
   52740: out<=0;
   52741: out<=1;
   52742: out<=0;
   52743: out<=1;
   52744: out<=1;
   52745: out<=0;
   52746: out<=0;
   52747: out<=1;
   52748: out<=0;
   52749: out<=0;
   52750: out<=0;
   52751: out<=0;
   52752: out<=1;
   52753: out<=0;
   52754: out<=1;
   52755: out<=0;
   52756: out<=1;
   52757: out<=1;
   52758: out<=0;
   52759: out<=0;
   52760: out<=0;
   52761: out<=0;
   52762: out<=0;
   52763: out<=0;
   52764: out<=0;
   52765: out<=1;
   52766: out<=1;
   52767: out<=0;
   52768: out<=1;
   52769: out<=0;
   52770: out<=0;
   52771: out<=1;
   52772: out<=1;
   52773: out<=1;
   52774: out<=1;
   52775: out<=1;
   52776: out<=1;
   52777: out<=1;
   52778: out<=0;
   52779: out<=0;
   52780: out<=1;
   52781: out<=0;
   52782: out<=1;
   52783: out<=0;
   52784: out<=1;
   52785: out<=1;
   52786: out<=1;
   52787: out<=1;
   52788: out<=0;
   52789: out<=1;
   52790: out<=1;
   52791: out<=0;
   52792: out<=0;
   52793: out<=1;
   52794: out<=0;
   52795: out<=1;
   52796: out<=1;
   52797: out<=1;
   52798: out<=0;
   52799: out<=0;
   52800: out<=1;
   52801: out<=1;
   52802: out<=0;
   52803: out<=0;
   52804: out<=0;
   52805: out<=1;
   52806: out<=0;
   52807: out<=1;
   52808: out<=1;
   52809: out<=0;
   52810: out<=0;
   52811: out<=1;
   52812: out<=0;
   52813: out<=0;
   52814: out<=0;
   52815: out<=0;
   52816: out<=0;
   52817: out<=1;
   52818: out<=0;
   52819: out<=1;
   52820: out<=0;
   52821: out<=0;
   52822: out<=1;
   52823: out<=1;
   52824: out<=1;
   52825: out<=1;
   52826: out<=1;
   52827: out<=1;
   52828: out<=1;
   52829: out<=0;
   52830: out<=0;
   52831: out<=1;
   52832: out<=0;
   52833: out<=1;
   52834: out<=1;
   52835: out<=0;
   52836: out<=0;
   52837: out<=0;
   52838: out<=0;
   52839: out<=0;
   52840: out<=0;
   52841: out<=0;
   52842: out<=1;
   52843: out<=1;
   52844: out<=0;
   52845: out<=1;
   52846: out<=0;
   52847: out<=1;
   52848: out<=1;
   52849: out<=1;
   52850: out<=1;
   52851: out<=1;
   52852: out<=0;
   52853: out<=1;
   52854: out<=1;
   52855: out<=0;
   52856: out<=0;
   52857: out<=1;
   52858: out<=0;
   52859: out<=1;
   52860: out<=1;
   52861: out<=1;
   52862: out<=0;
   52863: out<=0;
   52864: out<=1;
   52865: out<=1;
   52866: out<=0;
   52867: out<=0;
   52868: out<=0;
   52869: out<=1;
   52870: out<=0;
   52871: out<=1;
   52872: out<=1;
   52873: out<=0;
   52874: out<=0;
   52875: out<=1;
   52876: out<=0;
   52877: out<=0;
   52878: out<=0;
   52879: out<=0;
   52880: out<=0;
   52881: out<=1;
   52882: out<=0;
   52883: out<=1;
   52884: out<=0;
   52885: out<=0;
   52886: out<=1;
   52887: out<=1;
   52888: out<=1;
   52889: out<=1;
   52890: out<=1;
   52891: out<=1;
   52892: out<=1;
   52893: out<=0;
   52894: out<=0;
   52895: out<=1;
   52896: out<=1;
   52897: out<=0;
   52898: out<=0;
   52899: out<=1;
   52900: out<=1;
   52901: out<=1;
   52902: out<=1;
   52903: out<=1;
   52904: out<=1;
   52905: out<=1;
   52906: out<=0;
   52907: out<=0;
   52908: out<=1;
   52909: out<=0;
   52910: out<=1;
   52911: out<=0;
   52912: out<=0;
   52913: out<=0;
   52914: out<=0;
   52915: out<=0;
   52916: out<=1;
   52917: out<=0;
   52918: out<=0;
   52919: out<=1;
   52920: out<=1;
   52921: out<=0;
   52922: out<=1;
   52923: out<=0;
   52924: out<=0;
   52925: out<=0;
   52926: out<=1;
   52927: out<=1;
   52928: out<=1;
   52929: out<=1;
   52930: out<=0;
   52931: out<=0;
   52932: out<=0;
   52933: out<=1;
   52934: out<=0;
   52935: out<=1;
   52936: out<=1;
   52937: out<=0;
   52938: out<=0;
   52939: out<=1;
   52940: out<=0;
   52941: out<=0;
   52942: out<=0;
   52943: out<=0;
   52944: out<=1;
   52945: out<=0;
   52946: out<=1;
   52947: out<=0;
   52948: out<=1;
   52949: out<=1;
   52950: out<=0;
   52951: out<=0;
   52952: out<=0;
   52953: out<=0;
   52954: out<=0;
   52955: out<=0;
   52956: out<=0;
   52957: out<=1;
   52958: out<=1;
   52959: out<=0;
   52960: out<=0;
   52961: out<=1;
   52962: out<=1;
   52963: out<=0;
   52964: out<=0;
   52965: out<=0;
   52966: out<=0;
   52967: out<=0;
   52968: out<=0;
   52969: out<=0;
   52970: out<=1;
   52971: out<=1;
   52972: out<=0;
   52973: out<=1;
   52974: out<=0;
   52975: out<=1;
   52976: out<=0;
   52977: out<=0;
   52978: out<=0;
   52979: out<=0;
   52980: out<=1;
   52981: out<=0;
   52982: out<=0;
   52983: out<=1;
   52984: out<=1;
   52985: out<=0;
   52986: out<=1;
   52987: out<=0;
   52988: out<=0;
   52989: out<=0;
   52990: out<=1;
   52991: out<=1;
   52992: out<=0;
   52993: out<=1;
   52994: out<=0;
   52995: out<=1;
   52996: out<=0;
   52997: out<=0;
   52998: out<=1;
   52999: out<=1;
   53000: out<=1;
   53001: out<=1;
   53002: out<=1;
   53003: out<=1;
   53004: out<=1;
   53005: out<=0;
   53006: out<=0;
   53007: out<=1;
   53008: out<=1;
   53009: out<=1;
   53010: out<=0;
   53011: out<=0;
   53012: out<=0;
   53013: out<=1;
   53014: out<=0;
   53015: out<=1;
   53016: out<=1;
   53017: out<=0;
   53018: out<=0;
   53019: out<=1;
   53020: out<=0;
   53021: out<=0;
   53022: out<=0;
   53023: out<=0;
   53024: out<=1;
   53025: out<=1;
   53026: out<=1;
   53027: out<=1;
   53028: out<=0;
   53029: out<=1;
   53030: out<=1;
   53031: out<=0;
   53032: out<=0;
   53033: out<=1;
   53034: out<=0;
   53035: out<=1;
   53036: out<=1;
   53037: out<=1;
   53038: out<=0;
   53039: out<=0;
   53040: out<=0;
   53041: out<=1;
   53042: out<=1;
   53043: out<=0;
   53044: out<=0;
   53045: out<=0;
   53046: out<=0;
   53047: out<=0;
   53048: out<=0;
   53049: out<=0;
   53050: out<=1;
   53051: out<=1;
   53052: out<=0;
   53053: out<=1;
   53054: out<=0;
   53055: out<=1;
   53056: out<=1;
   53057: out<=0;
   53058: out<=1;
   53059: out<=0;
   53060: out<=1;
   53061: out<=1;
   53062: out<=0;
   53063: out<=0;
   53064: out<=0;
   53065: out<=0;
   53066: out<=0;
   53067: out<=0;
   53068: out<=0;
   53069: out<=1;
   53070: out<=1;
   53071: out<=0;
   53072: out<=1;
   53073: out<=1;
   53074: out<=0;
   53075: out<=0;
   53076: out<=0;
   53077: out<=1;
   53078: out<=0;
   53079: out<=1;
   53080: out<=1;
   53081: out<=0;
   53082: out<=0;
   53083: out<=1;
   53084: out<=0;
   53085: out<=0;
   53086: out<=0;
   53087: out<=0;
   53088: out<=1;
   53089: out<=1;
   53090: out<=1;
   53091: out<=1;
   53092: out<=0;
   53093: out<=1;
   53094: out<=1;
   53095: out<=0;
   53096: out<=0;
   53097: out<=1;
   53098: out<=0;
   53099: out<=1;
   53100: out<=1;
   53101: out<=1;
   53102: out<=0;
   53103: out<=0;
   53104: out<=1;
   53105: out<=0;
   53106: out<=0;
   53107: out<=1;
   53108: out<=1;
   53109: out<=1;
   53110: out<=1;
   53111: out<=1;
   53112: out<=1;
   53113: out<=1;
   53114: out<=0;
   53115: out<=0;
   53116: out<=1;
   53117: out<=0;
   53118: out<=1;
   53119: out<=0;
   53120: out<=1;
   53121: out<=0;
   53122: out<=1;
   53123: out<=0;
   53124: out<=1;
   53125: out<=1;
   53126: out<=0;
   53127: out<=0;
   53128: out<=0;
   53129: out<=0;
   53130: out<=0;
   53131: out<=0;
   53132: out<=0;
   53133: out<=1;
   53134: out<=1;
   53135: out<=0;
   53136: out<=1;
   53137: out<=1;
   53138: out<=0;
   53139: out<=0;
   53140: out<=0;
   53141: out<=1;
   53142: out<=0;
   53143: out<=1;
   53144: out<=1;
   53145: out<=0;
   53146: out<=0;
   53147: out<=1;
   53148: out<=0;
   53149: out<=0;
   53150: out<=0;
   53151: out<=0;
   53152: out<=0;
   53153: out<=0;
   53154: out<=0;
   53155: out<=0;
   53156: out<=1;
   53157: out<=0;
   53158: out<=0;
   53159: out<=1;
   53160: out<=1;
   53161: out<=0;
   53162: out<=1;
   53163: out<=0;
   53164: out<=0;
   53165: out<=0;
   53166: out<=1;
   53167: out<=1;
   53168: out<=0;
   53169: out<=1;
   53170: out<=1;
   53171: out<=0;
   53172: out<=0;
   53173: out<=0;
   53174: out<=0;
   53175: out<=0;
   53176: out<=0;
   53177: out<=0;
   53178: out<=1;
   53179: out<=1;
   53180: out<=0;
   53181: out<=1;
   53182: out<=0;
   53183: out<=1;
   53184: out<=0;
   53185: out<=1;
   53186: out<=0;
   53187: out<=1;
   53188: out<=0;
   53189: out<=0;
   53190: out<=1;
   53191: out<=1;
   53192: out<=1;
   53193: out<=1;
   53194: out<=1;
   53195: out<=1;
   53196: out<=1;
   53197: out<=0;
   53198: out<=0;
   53199: out<=1;
   53200: out<=1;
   53201: out<=1;
   53202: out<=0;
   53203: out<=0;
   53204: out<=0;
   53205: out<=1;
   53206: out<=0;
   53207: out<=1;
   53208: out<=1;
   53209: out<=0;
   53210: out<=0;
   53211: out<=1;
   53212: out<=0;
   53213: out<=0;
   53214: out<=0;
   53215: out<=0;
   53216: out<=0;
   53217: out<=0;
   53218: out<=0;
   53219: out<=0;
   53220: out<=1;
   53221: out<=0;
   53222: out<=0;
   53223: out<=1;
   53224: out<=1;
   53225: out<=0;
   53226: out<=1;
   53227: out<=0;
   53228: out<=0;
   53229: out<=0;
   53230: out<=1;
   53231: out<=1;
   53232: out<=1;
   53233: out<=0;
   53234: out<=0;
   53235: out<=1;
   53236: out<=1;
   53237: out<=1;
   53238: out<=1;
   53239: out<=1;
   53240: out<=1;
   53241: out<=1;
   53242: out<=0;
   53243: out<=0;
   53244: out<=1;
   53245: out<=0;
   53246: out<=1;
   53247: out<=0;
   53248: out<=0;
   53249: out<=1;
   53250: out<=0;
   53251: out<=1;
   53252: out<=1;
   53253: out<=1;
   53254: out<=0;
   53255: out<=0;
   53256: out<=1;
   53257: out<=1;
   53258: out<=1;
   53259: out<=1;
   53260: out<=0;
   53261: out<=1;
   53262: out<=1;
   53263: out<=0;
   53264: out<=1;
   53265: out<=1;
   53266: out<=0;
   53267: out<=0;
   53268: out<=1;
   53269: out<=0;
   53270: out<=1;
   53271: out<=0;
   53272: out<=1;
   53273: out<=0;
   53274: out<=0;
   53275: out<=1;
   53276: out<=1;
   53277: out<=1;
   53278: out<=1;
   53279: out<=1;
   53280: out<=0;
   53281: out<=0;
   53282: out<=0;
   53283: out<=0;
   53284: out<=0;
   53285: out<=1;
   53286: out<=1;
   53287: out<=0;
   53288: out<=1;
   53289: out<=0;
   53290: out<=1;
   53291: out<=0;
   53292: out<=1;
   53293: out<=1;
   53294: out<=0;
   53295: out<=0;
   53296: out<=1;
   53297: out<=0;
   53298: out<=0;
   53299: out<=1;
   53300: out<=0;
   53301: out<=0;
   53302: out<=0;
   53303: out<=0;
   53304: out<=1;
   53305: out<=1;
   53306: out<=0;
   53307: out<=0;
   53308: out<=0;
   53309: out<=1;
   53310: out<=0;
   53311: out<=1;
   53312: out<=1;
   53313: out<=0;
   53314: out<=1;
   53315: out<=0;
   53316: out<=0;
   53317: out<=0;
   53318: out<=1;
   53319: out<=1;
   53320: out<=0;
   53321: out<=0;
   53322: out<=0;
   53323: out<=0;
   53324: out<=1;
   53325: out<=0;
   53326: out<=0;
   53327: out<=1;
   53328: out<=1;
   53329: out<=1;
   53330: out<=0;
   53331: out<=0;
   53332: out<=1;
   53333: out<=0;
   53334: out<=1;
   53335: out<=0;
   53336: out<=1;
   53337: out<=0;
   53338: out<=0;
   53339: out<=1;
   53340: out<=1;
   53341: out<=1;
   53342: out<=1;
   53343: out<=1;
   53344: out<=0;
   53345: out<=0;
   53346: out<=0;
   53347: out<=0;
   53348: out<=0;
   53349: out<=1;
   53350: out<=1;
   53351: out<=0;
   53352: out<=1;
   53353: out<=0;
   53354: out<=1;
   53355: out<=0;
   53356: out<=1;
   53357: out<=1;
   53358: out<=0;
   53359: out<=0;
   53360: out<=0;
   53361: out<=1;
   53362: out<=1;
   53363: out<=0;
   53364: out<=1;
   53365: out<=1;
   53366: out<=1;
   53367: out<=1;
   53368: out<=0;
   53369: out<=0;
   53370: out<=1;
   53371: out<=1;
   53372: out<=1;
   53373: out<=0;
   53374: out<=1;
   53375: out<=0;
   53376: out<=1;
   53377: out<=0;
   53378: out<=1;
   53379: out<=0;
   53380: out<=0;
   53381: out<=0;
   53382: out<=1;
   53383: out<=1;
   53384: out<=0;
   53385: out<=0;
   53386: out<=0;
   53387: out<=0;
   53388: out<=1;
   53389: out<=0;
   53390: out<=0;
   53391: out<=1;
   53392: out<=1;
   53393: out<=1;
   53394: out<=0;
   53395: out<=0;
   53396: out<=1;
   53397: out<=0;
   53398: out<=1;
   53399: out<=0;
   53400: out<=1;
   53401: out<=0;
   53402: out<=0;
   53403: out<=1;
   53404: out<=1;
   53405: out<=1;
   53406: out<=1;
   53407: out<=1;
   53408: out<=1;
   53409: out<=1;
   53410: out<=1;
   53411: out<=1;
   53412: out<=1;
   53413: out<=0;
   53414: out<=0;
   53415: out<=1;
   53416: out<=0;
   53417: out<=1;
   53418: out<=0;
   53419: out<=1;
   53420: out<=0;
   53421: out<=0;
   53422: out<=1;
   53423: out<=1;
   53424: out<=1;
   53425: out<=0;
   53426: out<=0;
   53427: out<=1;
   53428: out<=0;
   53429: out<=0;
   53430: out<=0;
   53431: out<=0;
   53432: out<=1;
   53433: out<=1;
   53434: out<=0;
   53435: out<=0;
   53436: out<=0;
   53437: out<=1;
   53438: out<=0;
   53439: out<=1;
   53440: out<=0;
   53441: out<=1;
   53442: out<=0;
   53443: out<=1;
   53444: out<=1;
   53445: out<=1;
   53446: out<=0;
   53447: out<=0;
   53448: out<=1;
   53449: out<=1;
   53450: out<=1;
   53451: out<=1;
   53452: out<=0;
   53453: out<=1;
   53454: out<=1;
   53455: out<=0;
   53456: out<=1;
   53457: out<=1;
   53458: out<=0;
   53459: out<=0;
   53460: out<=1;
   53461: out<=0;
   53462: out<=1;
   53463: out<=0;
   53464: out<=1;
   53465: out<=0;
   53466: out<=0;
   53467: out<=1;
   53468: out<=1;
   53469: out<=1;
   53470: out<=1;
   53471: out<=1;
   53472: out<=1;
   53473: out<=1;
   53474: out<=1;
   53475: out<=1;
   53476: out<=1;
   53477: out<=0;
   53478: out<=0;
   53479: out<=1;
   53480: out<=0;
   53481: out<=1;
   53482: out<=0;
   53483: out<=1;
   53484: out<=0;
   53485: out<=0;
   53486: out<=1;
   53487: out<=1;
   53488: out<=0;
   53489: out<=1;
   53490: out<=1;
   53491: out<=0;
   53492: out<=1;
   53493: out<=1;
   53494: out<=1;
   53495: out<=1;
   53496: out<=0;
   53497: out<=0;
   53498: out<=1;
   53499: out<=1;
   53500: out<=1;
   53501: out<=0;
   53502: out<=1;
   53503: out<=0;
   53504: out<=1;
   53505: out<=1;
   53506: out<=0;
   53507: out<=0;
   53508: out<=1;
   53509: out<=0;
   53510: out<=1;
   53511: out<=0;
   53512: out<=1;
   53513: out<=0;
   53514: out<=0;
   53515: out<=1;
   53516: out<=1;
   53517: out<=1;
   53518: out<=1;
   53519: out<=1;
   53520: out<=1;
   53521: out<=0;
   53522: out<=1;
   53523: out<=0;
   53524: out<=0;
   53525: out<=0;
   53526: out<=1;
   53527: out<=1;
   53528: out<=0;
   53529: out<=0;
   53530: out<=0;
   53531: out<=0;
   53532: out<=1;
   53533: out<=0;
   53534: out<=0;
   53535: out<=1;
   53536: out<=0;
   53537: out<=1;
   53538: out<=1;
   53539: out<=0;
   53540: out<=1;
   53541: out<=1;
   53542: out<=1;
   53543: out<=1;
   53544: out<=0;
   53545: out<=0;
   53546: out<=1;
   53547: out<=1;
   53548: out<=1;
   53549: out<=0;
   53550: out<=1;
   53551: out<=0;
   53552: out<=0;
   53553: out<=0;
   53554: out<=0;
   53555: out<=0;
   53556: out<=0;
   53557: out<=1;
   53558: out<=1;
   53559: out<=0;
   53560: out<=1;
   53561: out<=0;
   53562: out<=1;
   53563: out<=0;
   53564: out<=1;
   53565: out<=1;
   53566: out<=0;
   53567: out<=0;
   53568: out<=1;
   53569: out<=1;
   53570: out<=0;
   53571: out<=0;
   53572: out<=1;
   53573: out<=0;
   53574: out<=1;
   53575: out<=0;
   53576: out<=1;
   53577: out<=0;
   53578: out<=0;
   53579: out<=1;
   53580: out<=1;
   53581: out<=1;
   53582: out<=1;
   53583: out<=1;
   53584: out<=0;
   53585: out<=1;
   53586: out<=0;
   53587: out<=1;
   53588: out<=1;
   53589: out<=1;
   53590: out<=0;
   53591: out<=0;
   53592: out<=1;
   53593: out<=1;
   53594: out<=1;
   53595: out<=1;
   53596: out<=0;
   53597: out<=1;
   53598: out<=1;
   53599: out<=0;
   53600: out<=1;
   53601: out<=0;
   53602: out<=0;
   53603: out<=1;
   53604: out<=0;
   53605: out<=0;
   53606: out<=0;
   53607: out<=0;
   53608: out<=1;
   53609: out<=1;
   53610: out<=0;
   53611: out<=0;
   53612: out<=0;
   53613: out<=1;
   53614: out<=0;
   53615: out<=1;
   53616: out<=0;
   53617: out<=0;
   53618: out<=0;
   53619: out<=0;
   53620: out<=0;
   53621: out<=1;
   53622: out<=1;
   53623: out<=0;
   53624: out<=1;
   53625: out<=0;
   53626: out<=1;
   53627: out<=0;
   53628: out<=1;
   53629: out<=1;
   53630: out<=0;
   53631: out<=0;
   53632: out<=1;
   53633: out<=1;
   53634: out<=0;
   53635: out<=0;
   53636: out<=1;
   53637: out<=0;
   53638: out<=1;
   53639: out<=0;
   53640: out<=1;
   53641: out<=0;
   53642: out<=0;
   53643: out<=1;
   53644: out<=1;
   53645: out<=1;
   53646: out<=1;
   53647: out<=1;
   53648: out<=0;
   53649: out<=1;
   53650: out<=0;
   53651: out<=1;
   53652: out<=1;
   53653: out<=1;
   53654: out<=0;
   53655: out<=0;
   53656: out<=1;
   53657: out<=1;
   53658: out<=1;
   53659: out<=1;
   53660: out<=0;
   53661: out<=1;
   53662: out<=1;
   53663: out<=0;
   53664: out<=0;
   53665: out<=1;
   53666: out<=1;
   53667: out<=0;
   53668: out<=1;
   53669: out<=1;
   53670: out<=1;
   53671: out<=1;
   53672: out<=0;
   53673: out<=0;
   53674: out<=1;
   53675: out<=1;
   53676: out<=1;
   53677: out<=0;
   53678: out<=1;
   53679: out<=0;
   53680: out<=1;
   53681: out<=1;
   53682: out<=1;
   53683: out<=1;
   53684: out<=1;
   53685: out<=0;
   53686: out<=0;
   53687: out<=1;
   53688: out<=0;
   53689: out<=1;
   53690: out<=0;
   53691: out<=1;
   53692: out<=0;
   53693: out<=0;
   53694: out<=1;
   53695: out<=1;
   53696: out<=1;
   53697: out<=1;
   53698: out<=0;
   53699: out<=0;
   53700: out<=1;
   53701: out<=0;
   53702: out<=1;
   53703: out<=0;
   53704: out<=1;
   53705: out<=0;
   53706: out<=0;
   53707: out<=1;
   53708: out<=1;
   53709: out<=1;
   53710: out<=1;
   53711: out<=1;
   53712: out<=1;
   53713: out<=0;
   53714: out<=1;
   53715: out<=0;
   53716: out<=0;
   53717: out<=0;
   53718: out<=1;
   53719: out<=1;
   53720: out<=0;
   53721: out<=0;
   53722: out<=0;
   53723: out<=0;
   53724: out<=1;
   53725: out<=0;
   53726: out<=0;
   53727: out<=1;
   53728: out<=1;
   53729: out<=0;
   53730: out<=0;
   53731: out<=1;
   53732: out<=0;
   53733: out<=0;
   53734: out<=0;
   53735: out<=0;
   53736: out<=1;
   53737: out<=1;
   53738: out<=0;
   53739: out<=0;
   53740: out<=0;
   53741: out<=1;
   53742: out<=0;
   53743: out<=1;
   53744: out<=1;
   53745: out<=1;
   53746: out<=1;
   53747: out<=1;
   53748: out<=1;
   53749: out<=0;
   53750: out<=0;
   53751: out<=1;
   53752: out<=0;
   53753: out<=1;
   53754: out<=0;
   53755: out<=1;
   53756: out<=0;
   53757: out<=0;
   53758: out<=1;
   53759: out<=1;
   53760: out<=1;
   53761: out<=1;
   53762: out<=1;
   53763: out<=1;
   53764: out<=1;
   53765: out<=0;
   53766: out<=0;
   53767: out<=1;
   53768: out<=0;
   53769: out<=1;
   53770: out<=0;
   53771: out<=1;
   53772: out<=0;
   53773: out<=0;
   53774: out<=1;
   53775: out<=1;
   53776: out<=1;
   53777: out<=0;
   53778: out<=0;
   53779: out<=1;
   53780: out<=0;
   53781: out<=0;
   53782: out<=0;
   53783: out<=0;
   53784: out<=1;
   53785: out<=1;
   53786: out<=0;
   53787: out<=0;
   53788: out<=0;
   53789: out<=1;
   53790: out<=0;
   53791: out<=1;
   53792: out<=1;
   53793: out<=0;
   53794: out<=1;
   53795: out<=0;
   53796: out<=0;
   53797: out<=0;
   53798: out<=1;
   53799: out<=1;
   53800: out<=0;
   53801: out<=0;
   53802: out<=0;
   53803: out<=0;
   53804: out<=1;
   53805: out<=0;
   53806: out<=0;
   53807: out<=1;
   53808: out<=1;
   53809: out<=1;
   53810: out<=0;
   53811: out<=0;
   53812: out<=1;
   53813: out<=0;
   53814: out<=1;
   53815: out<=0;
   53816: out<=1;
   53817: out<=0;
   53818: out<=0;
   53819: out<=1;
   53820: out<=1;
   53821: out<=1;
   53822: out<=1;
   53823: out<=1;
   53824: out<=1;
   53825: out<=1;
   53826: out<=1;
   53827: out<=1;
   53828: out<=1;
   53829: out<=0;
   53830: out<=0;
   53831: out<=1;
   53832: out<=0;
   53833: out<=1;
   53834: out<=0;
   53835: out<=1;
   53836: out<=0;
   53837: out<=0;
   53838: out<=1;
   53839: out<=1;
   53840: out<=0;
   53841: out<=1;
   53842: out<=1;
   53843: out<=0;
   53844: out<=1;
   53845: out<=1;
   53846: out<=1;
   53847: out<=1;
   53848: out<=0;
   53849: out<=0;
   53850: out<=1;
   53851: out<=1;
   53852: out<=1;
   53853: out<=0;
   53854: out<=1;
   53855: out<=0;
   53856: out<=0;
   53857: out<=1;
   53858: out<=0;
   53859: out<=1;
   53860: out<=1;
   53861: out<=1;
   53862: out<=0;
   53863: out<=0;
   53864: out<=1;
   53865: out<=1;
   53866: out<=1;
   53867: out<=1;
   53868: out<=0;
   53869: out<=1;
   53870: out<=1;
   53871: out<=0;
   53872: out<=1;
   53873: out<=1;
   53874: out<=0;
   53875: out<=0;
   53876: out<=1;
   53877: out<=0;
   53878: out<=1;
   53879: out<=0;
   53880: out<=1;
   53881: out<=0;
   53882: out<=0;
   53883: out<=1;
   53884: out<=1;
   53885: out<=1;
   53886: out<=1;
   53887: out<=1;
   53888: out<=0;
   53889: out<=0;
   53890: out<=0;
   53891: out<=0;
   53892: out<=0;
   53893: out<=1;
   53894: out<=1;
   53895: out<=0;
   53896: out<=1;
   53897: out<=0;
   53898: out<=1;
   53899: out<=0;
   53900: out<=1;
   53901: out<=1;
   53902: out<=0;
   53903: out<=0;
   53904: out<=1;
   53905: out<=0;
   53906: out<=0;
   53907: out<=1;
   53908: out<=0;
   53909: out<=0;
   53910: out<=0;
   53911: out<=0;
   53912: out<=1;
   53913: out<=1;
   53914: out<=0;
   53915: out<=0;
   53916: out<=0;
   53917: out<=1;
   53918: out<=0;
   53919: out<=1;
   53920: out<=0;
   53921: out<=1;
   53922: out<=0;
   53923: out<=1;
   53924: out<=1;
   53925: out<=1;
   53926: out<=0;
   53927: out<=0;
   53928: out<=1;
   53929: out<=1;
   53930: out<=1;
   53931: out<=1;
   53932: out<=0;
   53933: out<=1;
   53934: out<=1;
   53935: out<=0;
   53936: out<=1;
   53937: out<=1;
   53938: out<=0;
   53939: out<=0;
   53940: out<=1;
   53941: out<=0;
   53942: out<=1;
   53943: out<=0;
   53944: out<=1;
   53945: out<=0;
   53946: out<=0;
   53947: out<=1;
   53948: out<=1;
   53949: out<=1;
   53950: out<=1;
   53951: out<=1;
   53952: out<=0;
   53953: out<=0;
   53954: out<=0;
   53955: out<=0;
   53956: out<=0;
   53957: out<=1;
   53958: out<=1;
   53959: out<=0;
   53960: out<=1;
   53961: out<=0;
   53962: out<=1;
   53963: out<=0;
   53964: out<=1;
   53965: out<=1;
   53966: out<=0;
   53967: out<=0;
   53968: out<=0;
   53969: out<=1;
   53970: out<=1;
   53971: out<=0;
   53972: out<=1;
   53973: out<=1;
   53974: out<=1;
   53975: out<=1;
   53976: out<=0;
   53977: out<=0;
   53978: out<=1;
   53979: out<=1;
   53980: out<=1;
   53981: out<=0;
   53982: out<=1;
   53983: out<=0;
   53984: out<=1;
   53985: out<=0;
   53986: out<=1;
   53987: out<=0;
   53988: out<=0;
   53989: out<=0;
   53990: out<=1;
   53991: out<=1;
   53992: out<=0;
   53993: out<=0;
   53994: out<=0;
   53995: out<=0;
   53996: out<=1;
   53997: out<=0;
   53998: out<=0;
   53999: out<=1;
   54000: out<=1;
   54001: out<=1;
   54002: out<=0;
   54003: out<=0;
   54004: out<=1;
   54005: out<=0;
   54006: out<=1;
   54007: out<=0;
   54008: out<=1;
   54009: out<=0;
   54010: out<=0;
   54011: out<=1;
   54012: out<=1;
   54013: out<=1;
   54014: out<=1;
   54015: out<=1;
   54016: out<=0;
   54017: out<=1;
   54018: out<=1;
   54019: out<=0;
   54020: out<=1;
   54021: out<=1;
   54022: out<=1;
   54023: out<=1;
   54024: out<=0;
   54025: out<=0;
   54026: out<=1;
   54027: out<=1;
   54028: out<=1;
   54029: out<=0;
   54030: out<=1;
   54031: out<=0;
   54032: out<=1;
   54033: out<=1;
   54034: out<=1;
   54035: out<=1;
   54036: out<=1;
   54037: out<=0;
   54038: out<=0;
   54039: out<=1;
   54040: out<=0;
   54041: out<=1;
   54042: out<=0;
   54043: out<=1;
   54044: out<=0;
   54045: out<=0;
   54046: out<=1;
   54047: out<=1;
   54048: out<=1;
   54049: out<=1;
   54050: out<=0;
   54051: out<=0;
   54052: out<=1;
   54053: out<=0;
   54054: out<=1;
   54055: out<=0;
   54056: out<=1;
   54057: out<=0;
   54058: out<=0;
   54059: out<=1;
   54060: out<=1;
   54061: out<=1;
   54062: out<=1;
   54063: out<=1;
   54064: out<=0;
   54065: out<=1;
   54066: out<=0;
   54067: out<=1;
   54068: out<=1;
   54069: out<=1;
   54070: out<=0;
   54071: out<=0;
   54072: out<=1;
   54073: out<=1;
   54074: out<=1;
   54075: out<=1;
   54076: out<=0;
   54077: out<=1;
   54078: out<=1;
   54079: out<=0;
   54080: out<=1;
   54081: out<=0;
   54082: out<=0;
   54083: out<=1;
   54084: out<=0;
   54085: out<=0;
   54086: out<=0;
   54087: out<=0;
   54088: out<=1;
   54089: out<=1;
   54090: out<=0;
   54091: out<=0;
   54092: out<=0;
   54093: out<=1;
   54094: out<=0;
   54095: out<=1;
   54096: out<=1;
   54097: out<=1;
   54098: out<=1;
   54099: out<=1;
   54100: out<=1;
   54101: out<=0;
   54102: out<=0;
   54103: out<=1;
   54104: out<=0;
   54105: out<=1;
   54106: out<=0;
   54107: out<=1;
   54108: out<=0;
   54109: out<=0;
   54110: out<=1;
   54111: out<=1;
   54112: out<=1;
   54113: out<=1;
   54114: out<=0;
   54115: out<=0;
   54116: out<=1;
   54117: out<=0;
   54118: out<=1;
   54119: out<=0;
   54120: out<=1;
   54121: out<=0;
   54122: out<=0;
   54123: out<=1;
   54124: out<=1;
   54125: out<=1;
   54126: out<=1;
   54127: out<=1;
   54128: out<=1;
   54129: out<=0;
   54130: out<=1;
   54131: out<=0;
   54132: out<=0;
   54133: out<=0;
   54134: out<=1;
   54135: out<=1;
   54136: out<=0;
   54137: out<=0;
   54138: out<=0;
   54139: out<=0;
   54140: out<=1;
   54141: out<=0;
   54142: out<=0;
   54143: out<=1;
   54144: out<=0;
   54145: out<=1;
   54146: out<=1;
   54147: out<=0;
   54148: out<=1;
   54149: out<=1;
   54150: out<=1;
   54151: out<=1;
   54152: out<=0;
   54153: out<=0;
   54154: out<=1;
   54155: out<=1;
   54156: out<=1;
   54157: out<=0;
   54158: out<=1;
   54159: out<=0;
   54160: out<=0;
   54161: out<=0;
   54162: out<=0;
   54163: out<=0;
   54164: out<=0;
   54165: out<=1;
   54166: out<=1;
   54167: out<=0;
   54168: out<=1;
   54169: out<=0;
   54170: out<=1;
   54171: out<=0;
   54172: out<=1;
   54173: out<=1;
   54174: out<=0;
   54175: out<=0;
   54176: out<=1;
   54177: out<=1;
   54178: out<=0;
   54179: out<=0;
   54180: out<=1;
   54181: out<=0;
   54182: out<=1;
   54183: out<=0;
   54184: out<=1;
   54185: out<=0;
   54186: out<=0;
   54187: out<=1;
   54188: out<=1;
   54189: out<=1;
   54190: out<=1;
   54191: out<=1;
   54192: out<=1;
   54193: out<=0;
   54194: out<=1;
   54195: out<=0;
   54196: out<=0;
   54197: out<=0;
   54198: out<=1;
   54199: out<=1;
   54200: out<=0;
   54201: out<=0;
   54202: out<=0;
   54203: out<=0;
   54204: out<=1;
   54205: out<=0;
   54206: out<=0;
   54207: out<=1;
   54208: out<=1;
   54209: out<=0;
   54210: out<=0;
   54211: out<=1;
   54212: out<=0;
   54213: out<=0;
   54214: out<=0;
   54215: out<=0;
   54216: out<=1;
   54217: out<=1;
   54218: out<=0;
   54219: out<=0;
   54220: out<=0;
   54221: out<=1;
   54222: out<=0;
   54223: out<=1;
   54224: out<=0;
   54225: out<=0;
   54226: out<=0;
   54227: out<=0;
   54228: out<=0;
   54229: out<=1;
   54230: out<=1;
   54231: out<=0;
   54232: out<=1;
   54233: out<=0;
   54234: out<=1;
   54235: out<=0;
   54236: out<=1;
   54237: out<=1;
   54238: out<=0;
   54239: out<=0;
   54240: out<=1;
   54241: out<=1;
   54242: out<=0;
   54243: out<=0;
   54244: out<=1;
   54245: out<=0;
   54246: out<=1;
   54247: out<=0;
   54248: out<=1;
   54249: out<=0;
   54250: out<=0;
   54251: out<=1;
   54252: out<=1;
   54253: out<=1;
   54254: out<=1;
   54255: out<=1;
   54256: out<=0;
   54257: out<=1;
   54258: out<=0;
   54259: out<=1;
   54260: out<=1;
   54261: out<=1;
   54262: out<=0;
   54263: out<=0;
   54264: out<=1;
   54265: out<=1;
   54266: out<=1;
   54267: out<=1;
   54268: out<=0;
   54269: out<=1;
   54270: out<=1;
   54271: out<=0;
   54272: out<=1;
   54273: out<=1;
   54274: out<=0;
   54275: out<=0;
   54276: out<=0;
   54277: out<=1;
   54278: out<=0;
   54279: out<=1;
   54280: out<=0;
   54281: out<=1;
   54282: out<=1;
   54283: out<=0;
   54284: out<=1;
   54285: out<=1;
   54286: out<=1;
   54287: out<=1;
   54288: out<=0;
   54289: out<=1;
   54290: out<=0;
   54291: out<=1;
   54292: out<=0;
   54293: out<=0;
   54294: out<=1;
   54295: out<=1;
   54296: out<=0;
   54297: out<=0;
   54298: out<=0;
   54299: out<=0;
   54300: out<=0;
   54301: out<=1;
   54302: out<=1;
   54303: out<=0;
   54304: out<=1;
   54305: out<=0;
   54306: out<=0;
   54307: out<=1;
   54308: out<=1;
   54309: out<=1;
   54310: out<=1;
   54311: out<=1;
   54312: out<=0;
   54313: out<=0;
   54314: out<=1;
   54315: out<=1;
   54316: out<=0;
   54317: out<=1;
   54318: out<=0;
   54319: out<=1;
   54320: out<=0;
   54321: out<=0;
   54322: out<=0;
   54323: out<=0;
   54324: out<=1;
   54325: out<=0;
   54326: out<=0;
   54327: out<=1;
   54328: out<=0;
   54329: out<=1;
   54330: out<=0;
   54331: out<=1;
   54332: out<=1;
   54333: out<=1;
   54334: out<=0;
   54335: out<=0;
   54336: out<=1;
   54337: out<=1;
   54338: out<=0;
   54339: out<=0;
   54340: out<=0;
   54341: out<=1;
   54342: out<=0;
   54343: out<=1;
   54344: out<=0;
   54345: out<=1;
   54346: out<=1;
   54347: out<=0;
   54348: out<=1;
   54349: out<=1;
   54350: out<=1;
   54351: out<=1;
   54352: out<=1;
   54353: out<=0;
   54354: out<=1;
   54355: out<=0;
   54356: out<=1;
   54357: out<=1;
   54358: out<=0;
   54359: out<=0;
   54360: out<=1;
   54361: out<=1;
   54362: out<=1;
   54363: out<=1;
   54364: out<=1;
   54365: out<=0;
   54366: out<=0;
   54367: out<=1;
   54368: out<=0;
   54369: out<=1;
   54370: out<=1;
   54371: out<=0;
   54372: out<=0;
   54373: out<=0;
   54374: out<=0;
   54375: out<=0;
   54376: out<=1;
   54377: out<=1;
   54378: out<=0;
   54379: out<=0;
   54380: out<=1;
   54381: out<=0;
   54382: out<=1;
   54383: out<=0;
   54384: out<=0;
   54385: out<=0;
   54386: out<=0;
   54387: out<=0;
   54388: out<=1;
   54389: out<=0;
   54390: out<=0;
   54391: out<=1;
   54392: out<=0;
   54393: out<=1;
   54394: out<=0;
   54395: out<=1;
   54396: out<=1;
   54397: out<=1;
   54398: out<=0;
   54399: out<=0;
   54400: out<=1;
   54401: out<=1;
   54402: out<=0;
   54403: out<=0;
   54404: out<=0;
   54405: out<=1;
   54406: out<=0;
   54407: out<=1;
   54408: out<=0;
   54409: out<=1;
   54410: out<=1;
   54411: out<=0;
   54412: out<=1;
   54413: out<=1;
   54414: out<=1;
   54415: out<=1;
   54416: out<=1;
   54417: out<=0;
   54418: out<=1;
   54419: out<=0;
   54420: out<=1;
   54421: out<=1;
   54422: out<=0;
   54423: out<=0;
   54424: out<=1;
   54425: out<=1;
   54426: out<=1;
   54427: out<=1;
   54428: out<=1;
   54429: out<=0;
   54430: out<=0;
   54431: out<=1;
   54432: out<=1;
   54433: out<=0;
   54434: out<=0;
   54435: out<=1;
   54436: out<=1;
   54437: out<=1;
   54438: out<=1;
   54439: out<=1;
   54440: out<=0;
   54441: out<=0;
   54442: out<=1;
   54443: out<=1;
   54444: out<=0;
   54445: out<=1;
   54446: out<=0;
   54447: out<=1;
   54448: out<=1;
   54449: out<=1;
   54450: out<=1;
   54451: out<=1;
   54452: out<=0;
   54453: out<=1;
   54454: out<=1;
   54455: out<=0;
   54456: out<=1;
   54457: out<=0;
   54458: out<=1;
   54459: out<=0;
   54460: out<=0;
   54461: out<=0;
   54462: out<=1;
   54463: out<=1;
   54464: out<=1;
   54465: out<=1;
   54466: out<=0;
   54467: out<=0;
   54468: out<=0;
   54469: out<=1;
   54470: out<=0;
   54471: out<=1;
   54472: out<=0;
   54473: out<=1;
   54474: out<=1;
   54475: out<=0;
   54476: out<=1;
   54477: out<=1;
   54478: out<=1;
   54479: out<=1;
   54480: out<=0;
   54481: out<=1;
   54482: out<=0;
   54483: out<=1;
   54484: out<=0;
   54485: out<=0;
   54486: out<=1;
   54487: out<=1;
   54488: out<=0;
   54489: out<=0;
   54490: out<=0;
   54491: out<=0;
   54492: out<=0;
   54493: out<=1;
   54494: out<=1;
   54495: out<=0;
   54496: out<=0;
   54497: out<=1;
   54498: out<=1;
   54499: out<=0;
   54500: out<=0;
   54501: out<=0;
   54502: out<=0;
   54503: out<=0;
   54504: out<=1;
   54505: out<=1;
   54506: out<=0;
   54507: out<=0;
   54508: out<=1;
   54509: out<=0;
   54510: out<=1;
   54511: out<=0;
   54512: out<=1;
   54513: out<=1;
   54514: out<=1;
   54515: out<=1;
   54516: out<=0;
   54517: out<=1;
   54518: out<=1;
   54519: out<=0;
   54520: out<=1;
   54521: out<=0;
   54522: out<=1;
   54523: out<=0;
   54524: out<=0;
   54525: out<=0;
   54526: out<=1;
   54527: out<=1;
   54528: out<=1;
   54529: out<=0;
   54530: out<=1;
   54531: out<=0;
   54532: out<=1;
   54533: out<=1;
   54534: out<=0;
   54535: out<=0;
   54536: out<=1;
   54537: out<=1;
   54538: out<=1;
   54539: out<=1;
   54540: out<=1;
   54541: out<=0;
   54542: out<=0;
   54543: out<=1;
   54544: out<=1;
   54545: out<=1;
   54546: out<=0;
   54547: out<=0;
   54548: out<=0;
   54549: out<=1;
   54550: out<=0;
   54551: out<=1;
   54552: out<=0;
   54553: out<=1;
   54554: out<=1;
   54555: out<=0;
   54556: out<=1;
   54557: out<=1;
   54558: out<=1;
   54559: out<=1;
   54560: out<=0;
   54561: out<=0;
   54562: out<=0;
   54563: out<=0;
   54564: out<=1;
   54565: out<=0;
   54566: out<=0;
   54567: out<=1;
   54568: out<=0;
   54569: out<=1;
   54570: out<=0;
   54571: out<=1;
   54572: out<=1;
   54573: out<=1;
   54574: out<=0;
   54575: out<=0;
   54576: out<=0;
   54577: out<=1;
   54578: out<=1;
   54579: out<=0;
   54580: out<=0;
   54581: out<=0;
   54582: out<=0;
   54583: out<=0;
   54584: out<=1;
   54585: out<=1;
   54586: out<=0;
   54587: out<=0;
   54588: out<=1;
   54589: out<=0;
   54590: out<=1;
   54591: out<=0;
   54592: out<=0;
   54593: out<=1;
   54594: out<=0;
   54595: out<=1;
   54596: out<=0;
   54597: out<=0;
   54598: out<=1;
   54599: out<=1;
   54600: out<=0;
   54601: out<=0;
   54602: out<=0;
   54603: out<=0;
   54604: out<=0;
   54605: out<=1;
   54606: out<=1;
   54607: out<=0;
   54608: out<=1;
   54609: out<=1;
   54610: out<=0;
   54611: out<=0;
   54612: out<=0;
   54613: out<=1;
   54614: out<=0;
   54615: out<=1;
   54616: out<=0;
   54617: out<=1;
   54618: out<=1;
   54619: out<=0;
   54620: out<=1;
   54621: out<=1;
   54622: out<=1;
   54623: out<=1;
   54624: out<=0;
   54625: out<=0;
   54626: out<=0;
   54627: out<=0;
   54628: out<=1;
   54629: out<=0;
   54630: out<=0;
   54631: out<=1;
   54632: out<=0;
   54633: out<=1;
   54634: out<=0;
   54635: out<=1;
   54636: out<=1;
   54637: out<=1;
   54638: out<=0;
   54639: out<=0;
   54640: out<=1;
   54641: out<=0;
   54642: out<=0;
   54643: out<=1;
   54644: out<=1;
   54645: out<=1;
   54646: out<=1;
   54647: out<=1;
   54648: out<=0;
   54649: out<=0;
   54650: out<=1;
   54651: out<=1;
   54652: out<=0;
   54653: out<=1;
   54654: out<=0;
   54655: out<=1;
   54656: out<=0;
   54657: out<=1;
   54658: out<=0;
   54659: out<=1;
   54660: out<=0;
   54661: out<=0;
   54662: out<=1;
   54663: out<=1;
   54664: out<=0;
   54665: out<=0;
   54666: out<=0;
   54667: out<=0;
   54668: out<=0;
   54669: out<=1;
   54670: out<=1;
   54671: out<=0;
   54672: out<=1;
   54673: out<=1;
   54674: out<=0;
   54675: out<=0;
   54676: out<=0;
   54677: out<=1;
   54678: out<=0;
   54679: out<=1;
   54680: out<=0;
   54681: out<=1;
   54682: out<=1;
   54683: out<=0;
   54684: out<=1;
   54685: out<=1;
   54686: out<=1;
   54687: out<=1;
   54688: out<=1;
   54689: out<=1;
   54690: out<=1;
   54691: out<=1;
   54692: out<=0;
   54693: out<=1;
   54694: out<=1;
   54695: out<=0;
   54696: out<=1;
   54697: out<=0;
   54698: out<=1;
   54699: out<=0;
   54700: out<=0;
   54701: out<=0;
   54702: out<=1;
   54703: out<=1;
   54704: out<=0;
   54705: out<=1;
   54706: out<=1;
   54707: out<=0;
   54708: out<=0;
   54709: out<=0;
   54710: out<=0;
   54711: out<=0;
   54712: out<=1;
   54713: out<=1;
   54714: out<=0;
   54715: out<=0;
   54716: out<=1;
   54717: out<=0;
   54718: out<=1;
   54719: out<=0;
   54720: out<=1;
   54721: out<=0;
   54722: out<=1;
   54723: out<=0;
   54724: out<=1;
   54725: out<=1;
   54726: out<=0;
   54727: out<=0;
   54728: out<=1;
   54729: out<=1;
   54730: out<=1;
   54731: out<=1;
   54732: out<=1;
   54733: out<=0;
   54734: out<=0;
   54735: out<=1;
   54736: out<=1;
   54737: out<=1;
   54738: out<=0;
   54739: out<=0;
   54740: out<=0;
   54741: out<=1;
   54742: out<=0;
   54743: out<=1;
   54744: out<=0;
   54745: out<=1;
   54746: out<=1;
   54747: out<=0;
   54748: out<=1;
   54749: out<=1;
   54750: out<=1;
   54751: out<=1;
   54752: out<=1;
   54753: out<=1;
   54754: out<=1;
   54755: out<=1;
   54756: out<=0;
   54757: out<=1;
   54758: out<=1;
   54759: out<=0;
   54760: out<=1;
   54761: out<=0;
   54762: out<=1;
   54763: out<=0;
   54764: out<=0;
   54765: out<=0;
   54766: out<=1;
   54767: out<=1;
   54768: out<=1;
   54769: out<=0;
   54770: out<=0;
   54771: out<=1;
   54772: out<=1;
   54773: out<=1;
   54774: out<=1;
   54775: out<=1;
   54776: out<=0;
   54777: out<=0;
   54778: out<=1;
   54779: out<=1;
   54780: out<=0;
   54781: out<=1;
   54782: out<=0;
   54783: out<=1;
   54784: out<=1;
   54785: out<=0;
   54786: out<=0;
   54787: out<=1;
   54788: out<=1;
   54789: out<=1;
   54790: out<=1;
   54791: out<=1;
   54792: out<=0;
   54793: out<=0;
   54794: out<=1;
   54795: out<=1;
   54796: out<=0;
   54797: out<=1;
   54798: out<=0;
   54799: out<=1;
   54800: out<=1;
   54801: out<=1;
   54802: out<=1;
   54803: out<=1;
   54804: out<=0;
   54805: out<=1;
   54806: out<=1;
   54807: out<=0;
   54808: out<=1;
   54809: out<=0;
   54810: out<=1;
   54811: out<=0;
   54812: out<=0;
   54813: out<=0;
   54814: out<=1;
   54815: out<=1;
   54816: out<=1;
   54817: out<=1;
   54818: out<=0;
   54819: out<=0;
   54820: out<=0;
   54821: out<=1;
   54822: out<=0;
   54823: out<=1;
   54824: out<=0;
   54825: out<=1;
   54826: out<=1;
   54827: out<=0;
   54828: out<=1;
   54829: out<=1;
   54830: out<=1;
   54831: out<=1;
   54832: out<=1;
   54833: out<=0;
   54834: out<=1;
   54835: out<=0;
   54836: out<=1;
   54837: out<=1;
   54838: out<=0;
   54839: out<=0;
   54840: out<=1;
   54841: out<=1;
   54842: out<=1;
   54843: out<=1;
   54844: out<=1;
   54845: out<=0;
   54846: out<=0;
   54847: out<=1;
   54848: out<=0;
   54849: out<=1;
   54850: out<=1;
   54851: out<=0;
   54852: out<=0;
   54853: out<=0;
   54854: out<=0;
   54855: out<=0;
   54856: out<=1;
   54857: out<=1;
   54858: out<=0;
   54859: out<=0;
   54860: out<=1;
   54861: out<=0;
   54862: out<=1;
   54863: out<=0;
   54864: out<=1;
   54865: out<=1;
   54866: out<=1;
   54867: out<=1;
   54868: out<=0;
   54869: out<=1;
   54870: out<=1;
   54871: out<=0;
   54872: out<=1;
   54873: out<=0;
   54874: out<=1;
   54875: out<=0;
   54876: out<=0;
   54877: out<=0;
   54878: out<=1;
   54879: out<=1;
   54880: out<=1;
   54881: out<=1;
   54882: out<=0;
   54883: out<=0;
   54884: out<=0;
   54885: out<=1;
   54886: out<=0;
   54887: out<=1;
   54888: out<=0;
   54889: out<=1;
   54890: out<=1;
   54891: out<=0;
   54892: out<=1;
   54893: out<=1;
   54894: out<=1;
   54895: out<=1;
   54896: out<=0;
   54897: out<=1;
   54898: out<=0;
   54899: out<=1;
   54900: out<=0;
   54901: out<=0;
   54902: out<=1;
   54903: out<=1;
   54904: out<=0;
   54905: out<=0;
   54906: out<=0;
   54907: out<=0;
   54908: out<=0;
   54909: out<=1;
   54910: out<=1;
   54911: out<=0;
   54912: out<=1;
   54913: out<=0;
   54914: out<=0;
   54915: out<=1;
   54916: out<=1;
   54917: out<=1;
   54918: out<=1;
   54919: out<=1;
   54920: out<=0;
   54921: out<=0;
   54922: out<=1;
   54923: out<=1;
   54924: out<=0;
   54925: out<=1;
   54926: out<=0;
   54927: out<=1;
   54928: out<=0;
   54929: out<=0;
   54930: out<=0;
   54931: out<=0;
   54932: out<=1;
   54933: out<=0;
   54934: out<=0;
   54935: out<=1;
   54936: out<=0;
   54937: out<=1;
   54938: out<=0;
   54939: out<=1;
   54940: out<=1;
   54941: out<=1;
   54942: out<=0;
   54943: out<=0;
   54944: out<=1;
   54945: out<=1;
   54946: out<=0;
   54947: out<=0;
   54948: out<=0;
   54949: out<=1;
   54950: out<=0;
   54951: out<=1;
   54952: out<=0;
   54953: out<=1;
   54954: out<=1;
   54955: out<=0;
   54956: out<=1;
   54957: out<=1;
   54958: out<=1;
   54959: out<=1;
   54960: out<=0;
   54961: out<=1;
   54962: out<=0;
   54963: out<=1;
   54964: out<=0;
   54965: out<=0;
   54966: out<=1;
   54967: out<=1;
   54968: out<=0;
   54969: out<=0;
   54970: out<=0;
   54971: out<=0;
   54972: out<=0;
   54973: out<=1;
   54974: out<=1;
   54975: out<=0;
   54976: out<=0;
   54977: out<=1;
   54978: out<=1;
   54979: out<=0;
   54980: out<=0;
   54981: out<=0;
   54982: out<=0;
   54983: out<=0;
   54984: out<=1;
   54985: out<=1;
   54986: out<=0;
   54987: out<=0;
   54988: out<=1;
   54989: out<=0;
   54990: out<=1;
   54991: out<=0;
   54992: out<=0;
   54993: out<=0;
   54994: out<=0;
   54995: out<=0;
   54996: out<=1;
   54997: out<=0;
   54998: out<=0;
   54999: out<=1;
   55000: out<=0;
   55001: out<=1;
   55002: out<=0;
   55003: out<=1;
   55004: out<=1;
   55005: out<=1;
   55006: out<=0;
   55007: out<=0;
   55008: out<=1;
   55009: out<=1;
   55010: out<=0;
   55011: out<=0;
   55012: out<=0;
   55013: out<=1;
   55014: out<=0;
   55015: out<=1;
   55016: out<=0;
   55017: out<=1;
   55018: out<=1;
   55019: out<=0;
   55020: out<=1;
   55021: out<=1;
   55022: out<=1;
   55023: out<=1;
   55024: out<=1;
   55025: out<=0;
   55026: out<=1;
   55027: out<=0;
   55028: out<=1;
   55029: out<=1;
   55030: out<=0;
   55031: out<=0;
   55032: out<=1;
   55033: out<=1;
   55034: out<=1;
   55035: out<=1;
   55036: out<=1;
   55037: out<=0;
   55038: out<=0;
   55039: out<=1;
   55040: out<=1;
   55041: out<=1;
   55042: out<=1;
   55043: out<=1;
   55044: out<=0;
   55045: out<=1;
   55046: out<=1;
   55047: out<=0;
   55048: out<=1;
   55049: out<=0;
   55050: out<=1;
   55051: out<=0;
   55052: out<=0;
   55053: out<=0;
   55054: out<=1;
   55055: out<=1;
   55056: out<=0;
   55057: out<=1;
   55058: out<=1;
   55059: out<=0;
   55060: out<=0;
   55061: out<=0;
   55062: out<=0;
   55063: out<=0;
   55064: out<=1;
   55065: out<=1;
   55066: out<=0;
   55067: out<=0;
   55068: out<=1;
   55069: out<=0;
   55070: out<=1;
   55071: out<=0;
   55072: out<=0;
   55073: out<=1;
   55074: out<=0;
   55075: out<=1;
   55076: out<=0;
   55077: out<=0;
   55078: out<=1;
   55079: out<=1;
   55080: out<=0;
   55081: out<=0;
   55082: out<=0;
   55083: out<=0;
   55084: out<=0;
   55085: out<=1;
   55086: out<=1;
   55087: out<=0;
   55088: out<=1;
   55089: out<=1;
   55090: out<=0;
   55091: out<=0;
   55092: out<=0;
   55093: out<=1;
   55094: out<=0;
   55095: out<=1;
   55096: out<=0;
   55097: out<=1;
   55098: out<=1;
   55099: out<=0;
   55100: out<=1;
   55101: out<=1;
   55102: out<=1;
   55103: out<=1;
   55104: out<=1;
   55105: out<=1;
   55106: out<=1;
   55107: out<=1;
   55108: out<=0;
   55109: out<=1;
   55110: out<=1;
   55111: out<=0;
   55112: out<=1;
   55113: out<=0;
   55114: out<=1;
   55115: out<=0;
   55116: out<=0;
   55117: out<=0;
   55118: out<=1;
   55119: out<=1;
   55120: out<=1;
   55121: out<=0;
   55122: out<=0;
   55123: out<=1;
   55124: out<=1;
   55125: out<=1;
   55126: out<=1;
   55127: out<=1;
   55128: out<=0;
   55129: out<=0;
   55130: out<=1;
   55131: out<=1;
   55132: out<=0;
   55133: out<=1;
   55134: out<=0;
   55135: out<=1;
   55136: out<=1;
   55137: out<=0;
   55138: out<=1;
   55139: out<=0;
   55140: out<=1;
   55141: out<=1;
   55142: out<=0;
   55143: out<=0;
   55144: out<=1;
   55145: out<=1;
   55146: out<=1;
   55147: out<=1;
   55148: out<=1;
   55149: out<=0;
   55150: out<=0;
   55151: out<=1;
   55152: out<=1;
   55153: out<=1;
   55154: out<=0;
   55155: out<=0;
   55156: out<=0;
   55157: out<=1;
   55158: out<=0;
   55159: out<=1;
   55160: out<=0;
   55161: out<=1;
   55162: out<=1;
   55163: out<=0;
   55164: out<=1;
   55165: out<=1;
   55166: out<=1;
   55167: out<=1;
   55168: out<=0;
   55169: out<=0;
   55170: out<=0;
   55171: out<=0;
   55172: out<=1;
   55173: out<=0;
   55174: out<=0;
   55175: out<=1;
   55176: out<=0;
   55177: out<=1;
   55178: out<=0;
   55179: out<=1;
   55180: out<=1;
   55181: out<=1;
   55182: out<=0;
   55183: out<=0;
   55184: out<=0;
   55185: out<=1;
   55186: out<=1;
   55187: out<=0;
   55188: out<=0;
   55189: out<=0;
   55190: out<=0;
   55191: out<=0;
   55192: out<=1;
   55193: out<=1;
   55194: out<=0;
   55195: out<=0;
   55196: out<=1;
   55197: out<=0;
   55198: out<=1;
   55199: out<=0;
   55200: out<=1;
   55201: out<=0;
   55202: out<=1;
   55203: out<=0;
   55204: out<=1;
   55205: out<=1;
   55206: out<=0;
   55207: out<=0;
   55208: out<=1;
   55209: out<=1;
   55210: out<=1;
   55211: out<=1;
   55212: out<=1;
   55213: out<=0;
   55214: out<=0;
   55215: out<=1;
   55216: out<=1;
   55217: out<=1;
   55218: out<=0;
   55219: out<=0;
   55220: out<=0;
   55221: out<=1;
   55222: out<=0;
   55223: out<=1;
   55224: out<=0;
   55225: out<=1;
   55226: out<=1;
   55227: out<=0;
   55228: out<=1;
   55229: out<=1;
   55230: out<=1;
   55231: out<=1;
   55232: out<=0;
   55233: out<=0;
   55234: out<=0;
   55235: out<=0;
   55236: out<=1;
   55237: out<=0;
   55238: out<=0;
   55239: out<=1;
   55240: out<=0;
   55241: out<=1;
   55242: out<=0;
   55243: out<=1;
   55244: out<=1;
   55245: out<=1;
   55246: out<=0;
   55247: out<=0;
   55248: out<=1;
   55249: out<=0;
   55250: out<=0;
   55251: out<=1;
   55252: out<=1;
   55253: out<=1;
   55254: out<=1;
   55255: out<=1;
   55256: out<=0;
   55257: out<=0;
   55258: out<=1;
   55259: out<=1;
   55260: out<=0;
   55261: out<=1;
   55262: out<=0;
   55263: out<=1;
   55264: out<=0;
   55265: out<=1;
   55266: out<=0;
   55267: out<=1;
   55268: out<=0;
   55269: out<=0;
   55270: out<=1;
   55271: out<=1;
   55272: out<=0;
   55273: out<=0;
   55274: out<=0;
   55275: out<=0;
   55276: out<=0;
   55277: out<=1;
   55278: out<=1;
   55279: out<=0;
   55280: out<=1;
   55281: out<=1;
   55282: out<=0;
   55283: out<=0;
   55284: out<=0;
   55285: out<=1;
   55286: out<=0;
   55287: out<=1;
   55288: out<=0;
   55289: out<=1;
   55290: out<=1;
   55291: out<=0;
   55292: out<=1;
   55293: out<=1;
   55294: out<=1;
   55295: out<=1;
   55296: out<=1;
   55297: out<=1;
   55298: out<=1;
   55299: out<=1;
   55300: out<=0;
   55301: out<=1;
   55302: out<=1;
   55303: out<=0;
   55304: out<=0;
   55305: out<=1;
   55306: out<=0;
   55307: out<=1;
   55308: out<=1;
   55309: out<=1;
   55310: out<=0;
   55311: out<=0;
   55312: out<=0;
   55313: out<=1;
   55314: out<=1;
   55315: out<=0;
   55316: out<=0;
   55317: out<=0;
   55318: out<=0;
   55319: out<=0;
   55320: out<=0;
   55321: out<=0;
   55322: out<=1;
   55323: out<=1;
   55324: out<=0;
   55325: out<=1;
   55326: out<=0;
   55327: out<=1;
   55328: out<=1;
   55329: out<=0;
   55330: out<=1;
   55331: out<=0;
   55332: out<=1;
   55333: out<=1;
   55334: out<=0;
   55335: out<=0;
   55336: out<=0;
   55337: out<=0;
   55338: out<=0;
   55339: out<=0;
   55340: out<=0;
   55341: out<=1;
   55342: out<=1;
   55343: out<=0;
   55344: out<=0;
   55345: out<=0;
   55346: out<=1;
   55347: out<=1;
   55348: out<=1;
   55349: out<=0;
   55350: out<=1;
   55351: out<=0;
   55352: out<=0;
   55353: out<=1;
   55354: out<=1;
   55355: out<=0;
   55356: out<=1;
   55357: out<=1;
   55358: out<=1;
   55359: out<=1;
   55360: out<=1;
   55361: out<=1;
   55362: out<=1;
   55363: out<=1;
   55364: out<=0;
   55365: out<=1;
   55366: out<=1;
   55367: out<=0;
   55368: out<=0;
   55369: out<=1;
   55370: out<=0;
   55371: out<=1;
   55372: out<=1;
   55373: out<=1;
   55374: out<=0;
   55375: out<=0;
   55376: out<=1;
   55377: out<=0;
   55378: out<=0;
   55379: out<=1;
   55380: out<=1;
   55381: out<=1;
   55382: out<=1;
   55383: out<=1;
   55384: out<=1;
   55385: out<=1;
   55386: out<=0;
   55387: out<=0;
   55388: out<=1;
   55389: out<=0;
   55390: out<=1;
   55391: out<=0;
   55392: out<=0;
   55393: out<=1;
   55394: out<=0;
   55395: out<=1;
   55396: out<=0;
   55397: out<=0;
   55398: out<=1;
   55399: out<=1;
   55400: out<=1;
   55401: out<=1;
   55402: out<=1;
   55403: out<=1;
   55404: out<=1;
   55405: out<=0;
   55406: out<=0;
   55407: out<=1;
   55408: out<=0;
   55409: out<=0;
   55410: out<=1;
   55411: out<=1;
   55412: out<=1;
   55413: out<=0;
   55414: out<=1;
   55415: out<=0;
   55416: out<=0;
   55417: out<=1;
   55418: out<=1;
   55419: out<=0;
   55420: out<=1;
   55421: out<=1;
   55422: out<=1;
   55423: out<=1;
   55424: out<=0;
   55425: out<=0;
   55426: out<=0;
   55427: out<=0;
   55428: out<=1;
   55429: out<=0;
   55430: out<=0;
   55431: out<=1;
   55432: out<=1;
   55433: out<=0;
   55434: out<=1;
   55435: out<=0;
   55436: out<=0;
   55437: out<=0;
   55438: out<=1;
   55439: out<=1;
   55440: out<=0;
   55441: out<=1;
   55442: out<=1;
   55443: out<=0;
   55444: out<=0;
   55445: out<=0;
   55446: out<=0;
   55447: out<=0;
   55448: out<=0;
   55449: out<=0;
   55450: out<=1;
   55451: out<=1;
   55452: out<=0;
   55453: out<=1;
   55454: out<=0;
   55455: out<=1;
   55456: out<=0;
   55457: out<=1;
   55458: out<=0;
   55459: out<=1;
   55460: out<=0;
   55461: out<=0;
   55462: out<=1;
   55463: out<=1;
   55464: out<=1;
   55465: out<=1;
   55466: out<=1;
   55467: out<=1;
   55468: out<=1;
   55469: out<=0;
   55470: out<=0;
   55471: out<=1;
   55472: out<=0;
   55473: out<=0;
   55474: out<=1;
   55475: out<=1;
   55476: out<=1;
   55477: out<=0;
   55478: out<=1;
   55479: out<=0;
   55480: out<=0;
   55481: out<=1;
   55482: out<=1;
   55483: out<=0;
   55484: out<=1;
   55485: out<=1;
   55486: out<=1;
   55487: out<=1;
   55488: out<=0;
   55489: out<=0;
   55490: out<=0;
   55491: out<=0;
   55492: out<=1;
   55493: out<=0;
   55494: out<=0;
   55495: out<=1;
   55496: out<=1;
   55497: out<=0;
   55498: out<=1;
   55499: out<=0;
   55500: out<=0;
   55501: out<=0;
   55502: out<=1;
   55503: out<=1;
   55504: out<=1;
   55505: out<=0;
   55506: out<=0;
   55507: out<=1;
   55508: out<=1;
   55509: out<=1;
   55510: out<=1;
   55511: out<=1;
   55512: out<=1;
   55513: out<=1;
   55514: out<=0;
   55515: out<=0;
   55516: out<=1;
   55517: out<=0;
   55518: out<=1;
   55519: out<=0;
   55520: out<=1;
   55521: out<=0;
   55522: out<=1;
   55523: out<=0;
   55524: out<=1;
   55525: out<=1;
   55526: out<=0;
   55527: out<=0;
   55528: out<=0;
   55529: out<=0;
   55530: out<=0;
   55531: out<=0;
   55532: out<=0;
   55533: out<=1;
   55534: out<=1;
   55535: out<=0;
   55536: out<=0;
   55537: out<=0;
   55538: out<=1;
   55539: out<=1;
   55540: out<=1;
   55541: out<=0;
   55542: out<=1;
   55543: out<=0;
   55544: out<=0;
   55545: out<=1;
   55546: out<=1;
   55547: out<=0;
   55548: out<=1;
   55549: out<=1;
   55550: out<=1;
   55551: out<=1;
   55552: out<=1;
   55553: out<=0;
   55554: out<=0;
   55555: out<=1;
   55556: out<=1;
   55557: out<=1;
   55558: out<=1;
   55559: out<=1;
   55560: out<=1;
   55561: out<=1;
   55562: out<=0;
   55563: out<=0;
   55564: out<=1;
   55565: out<=0;
   55566: out<=1;
   55567: out<=0;
   55568: out<=1;
   55569: out<=1;
   55570: out<=1;
   55571: out<=1;
   55572: out<=0;
   55573: out<=1;
   55574: out<=1;
   55575: out<=0;
   55576: out<=0;
   55577: out<=1;
   55578: out<=0;
   55579: out<=1;
   55580: out<=1;
   55581: out<=1;
   55582: out<=0;
   55583: out<=0;
   55584: out<=0;
   55585: out<=0;
   55586: out<=1;
   55587: out<=1;
   55588: out<=1;
   55589: out<=0;
   55590: out<=1;
   55591: out<=0;
   55592: out<=0;
   55593: out<=1;
   55594: out<=1;
   55595: out<=0;
   55596: out<=1;
   55597: out<=1;
   55598: out<=1;
   55599: out<=1;
   55600: out<=0;
   55601: out<=1;
   55602: out<=0;
   55603: out<=1;
   55604: out<=0;
   55605: out<=0;
   55606: out<=1;
   55607: out<=1;
   55608: out<=1;
   55609: out<=1;
   55610: out<=1;
   55611: out<=1;
   55612: out<=1;
   55613: out<=0;
   55614: out<=0;
   55615: out<=1;
   55616: out<=0;
   55617: out<=1;
   55618: out<=1;
   55619: out<=0;
   55620: out<=0;
   55621: out<=0;
   55622: out<=0;
   55623: out<=0;
   55624: out<=0;
   55625: out<=0;
   55626: out<=1;
   55627: out<=1;
   55628: out<=0;
   55629: out<=1;
   55630: out<=0;
   55631: out<=1;
   55632: out<=1;
   55633: out<=1;
   55634: out<=1;
   55635: out<=1;
   55636: out<=0;
   55637: out<=1;
   55638: out<=1;
   55639: out<=0;
   55640: out<=0;
   55641: out<=1;
   55642: out<=0;
   55643: out<=1;
   55644: out<=1;
   55645: out<=1;
   55646: out<=0;
   55647: out<=0;
   55648: out<=0;
   55649: out<=0;
   55650: out<=1;
   55651: out<=1;
   55652: out<=1;
   55653: out<=0;
   55654: out<=1;
   55655: out<=0;
   55656: out<=0;
   55657: out<=1;
   55658: out<=1;
   55659: out<=0;
   55660: out<=1;
   55661: out<=1;
   55662: out<=1;
   55663: out<=1;
   55664: out<=1;
   55665: out<=0;
   55666: out<=1;
   55667: out<=0;
   55668: out<=1;
   55669: out<=1;
   55670: out<=0;
   55671: out<=0;
   55672: out<=0;
   55673: out<=0;
   55674: out<=0;
   55675: out<=0;
   55676: out<=0;
   55677: out<=1;
   55678: out<=1;
   55679: out<=0;
   55680: out<=1;
   55681: out<=0;
   55682: out<=0;
   55683: out<=1;
   55684: out<=1;
   55685: out<=1;
   55686: out<=1;
   55687: out<=1;
   55688: out<=1;
   55689: out<=1;
   55690: out<=0;
   55691: out<=0;
   55692: out<=1;
   55693: out<=0;
   55694: out<=1;
   55695: out<=0;
   55696: out<=0;
   55697: out<=0;
   55698: out<=0;
   55699: out<=0;
   55700: out<=1;
   55701: out<=0;
   55702: out<=0;
   55703: out<=1;
   55704: out<=1;
   55705: out<=0;
   55706: out<=1;
   55707: out<=0;
   55708: out<=0;
   55709: out<=0;
   55710: out<=1;
   55711: out<=1;
   55712: out<=0;
   55713: out<=0;
   55714: out<=1;
   55715: out<=1;
   55716: out<=1;
   55717: out<=0;
   55718: out<=1;
   55719: out<=0;
   55720: out<=0;
   55721: out<=1;
   55722: out<=1;
   55723: out<=0;
   55724: out<=1;
   55725: out<=1;
   55726: out<=1;
   55727: out<=1;
   55728: out<=1;
   55729: out<=0;
   55730: out<=1;
   55731: out<=0;
   55732: out<=1;
   55733: out<=1;
   55734: out<=0;
   55735: out<=0;
   55736: out<=0;
   55737: out<=0;
   55738: out<=0;
   55739: out<=0;
   55740: out<=0;
   55741: out<=1;
   55742: out<=1;
   55743: out<=0;
   55744: out<=0;
   55745: out<=1;
   55746: out<=1;
   55747: out<=0;
   55748: out<=0;
   55749: out<=0;
   55750: out<=0;
   55751: out<=0;
   55752: out<=0;
   55753: out<=0;
   55754: out<=1;
   55755: out<=1;
   55756: out<=0;
   55757: out<=1;
   55758: out<=0;
   55759: out<=1;
   55760: out<=0;
   55761: out<=0;
   55762: out<=0;
   55763: out<=0;
   55764: out<=1;
   55765: out<=0;
   55766: out<=0;
   55767: out<=1;
   55768: out<=1;
   55769: out<=0;
   55770: out<=1;
   55771: out<=0;
   55772: out<=0;
   55773: out<=0;
   55774: out<=1;
   55775: out<=1;
   55776: out<=0;
   55777: out<=0;
   55778: out<=1;
   55779: out<=1;
   55780: out<=1;
   55781: out<=0;
   55782: out<=1;
   55783: out<=0;
   55784: out<=0;
   55785: out<=1;
   55786: out<=1;
   55787: out<=0;
   55788: out<=1;
   55789: out<=1;
   55790: out<=1;
   55791: out<=1;
   55792: out<=0;
   55793: out<=1;
   55794: out<=0;
   55795: out<=1;
   55796: out<=0;
   55797: out<=0;
   55798: out<=1;
   55799: out<=1;
   55800: out<=1;
   55801: out<=1;
   55802: out<=1;
   55803: out<=1;
   55804: out<=1;
   55805: out<=0;
   55806: out<=0;
   55807: out<=1;
   55808: out<=0;
   55809: out<=1;
   55810: out<=0;
   55811: out<=1;
   55812: out<=0;
   55813: out<=0;
   55814: out<=1;
   55815: out<=1;
   55816: out<=1;
   55817: out<=1;
   55818: out<=1;
   55819: out<=1;
   55820: out<=1;
   55821: out<=0;
   55822: out<=0;
   55823: out<=1;
   55824: out<=0;
   55825: out<=0;
   55826: out<=1;
   55827: out<=1;
   55828: out<=1;
   55829: out<=0;
   55830: out<=1;
   55831: out<=0;
   55832: out<=0;
   55833: out<=1;
   55834: out<=1;
   55835: out<=0;
   55836: out<=1;
   55837: out<=1;
   55838: out<=1;
   55839: out<=1;
   55840: out<=0;
   55841: out<=0;
   55842: out<=0;
   55843: out<=0;
   55844: out<=1;
   55845: out<=0;
   55846: out<=0;
   55847: out<=1;
   55848: out<=1;
   55849: out<=0;
   55850: out<=1;
   55851: out<=0;
   55852: out<=0;
   55853: out<=0;
   55854: out<=1;
   55855: out<=1;
   55856: out<=0;
   55857: out<=1;
   55858: out<=1;
   55859: out<=0;
   55860: out<=0;
   55861: out<=0;
   55862: out<=0;
   55863: out<=0;
   55864: out<=0;
   55865: out<=0;
   55866: out<=1;
   55867: out<=1;
   55868: out<=0;
   55869: out<=1;
   55870: out<=0;
   55871: out<=1;
   55872: out<=1;
   55873: out<=0;
   55874: out<=1;
   55875: out<=0;
   55876: out<=1;
   55877: out<=1;
   55878: out<=0;
   55879: out<=0;
   55880: out<=0;
   55881: out<=0;
   55882: out<=0;
   55883: out<=0;
   55884: out<=0;
   55885: out<=1;
   55886: out<=1;
   55887: out<=0;
   55888: out<=0;
   55889: out<=0;
   55890: out<=1;
   55891: out<=1;
   55892: out<=1;
   55893: out<=0;
   55894: out<=1;
   55895: out<=0;
   55896: out<=0;
   55897: out<=1;
   55898: out<=1;
   55899: out<=0;
   55900: out<=1;
   55901: out<=1;
   55902: out<=1;
   55903: out<=1;
   55904: out<=0;
   55905: out<=0;
   55906: out<=0;
   55907: out<=0;
   55908: out<=1;
   55909: out<=0;
   55910: out<=0;
   55911: out<=1;
   55912: out<=1;
   55913: out<=0;
   55914: out<=1;
   55915: out<=0;
   55916: out<=0;
   55917: out<=0;
   55918: out<=1;
   55919: out<=1;
   55920: out<=1;
   55921: out<=0;
   55922: out<=0;
   55923: out<=1;
   55924: out<=1;
   55925: out<=1;
   55926: out<=1;
   55927: out<=1;
   55928: out<=1;
   55929: out<=1;
   55930: out<=0;
   55931: out<=0;
   55932: out<=1;
   55933: out<=0;
   55934: out<=1;
   55935: out<=0;
   55936: out<=1;
   55937: out<=0;
   55938: out<=1;
   55939: out<=0;
   55940: out<=1;
   55941: out<=1;
   55942: out<=0;
   55943: out<=0;
   55944: out<=0;
   55945: out<=0;
   55946: out<=0;
   55947: out<=0;
   55948: out<=0;
   55949: out<=1;
   55950: out<=1;
   55951: out<=0;
   55952: out<=0;
   55953: out<=0;
   55954: out<=1;
   55955: out<=1;
   55956: out<=1;
   55957: out<=0;
   55958: out<=1;
   55959: out<=0;
   55960: out<=0;
   55961: out<=1;
   55962: out<=1;
   55963: out<=0;
   55964: out<=1;
   55965: out<=1;
   55966: out<=1;
   55967: out<=1;
   55968: out<=1;
   55969: out<=1;
   55970: out<=1;
   55971: out<=1;
   55972: out<=0;
   55973: out<=1;
   55974: out<=1;
   55975: out<=0;
   55976: out<=0;
   55977: out<=1;
   55978: out<=0;
   55979: out<=1;
   55980: out<=1;
   55981: out<=1;
   55982: out<=0;
   55983: out<=0;
   55984: out<=0;
   55985: out<=1;
   55986: out<=1;
   55987: out<=0;
   55988: out<=0;
   55989: out<=0;
   55990: out<=0;
   55991: out<=0;
   55992: out<=0;
   55993: out<=0;
   55994: out<=1;
   55995: out<=1;
   55996: out<=0;
   55997: out<=1;
   55998: out<=0;
   55999: out<=1;
   56000: out<=0;
   56001: out<=1;
   56002: out<=0;
   56003: out<=1;
   56004: out<=0;
   56005: out<=0;
   56006: out<=1;
   56007: out<=1;
   56008: out<=1;
   56009: out<=1;
   56010: out<=1;
   56011: out<=1;
   56012: out<=1;
   56013: out<=0;
   56014: out<=0;
   56015: out<=1;
   56016: out<=0;
   56017: out<=0;
   56018: out<=1;
   56019: out<=1;
   56020: out<=1;
   56021: out<=0;
   56022: out<=1;
   56023: out<=0;
   56024: out<=0;
   56025: out<=1;
   56026: out<=1;
   56027: out<=0;
   56028: out<=1;
   56029: out<=1;
   56030: out<=1;
   56031: out<=1;
   56032: out<=1;
   56033: out<=1;
   56034: out<=1;
   56035: out<=1;
   56036: out<=0;
   56037: out<=1;
   56038: out<=1;
   56039: out<=0;
   56040: out<=0;
   56041: out<=1;
   56042: out<=0;
   56043: out<=1;
   56044: out<=1;
   56045: out<=1;
   56046: out<=0;
   56047: out<=0;
   56048: out<=1;
   56049: out<=0;
   56050: out<=0;
   56051: out<=1;
   56052: out<=1;
   56053: out<=1;
   56054: out<=1;
   56055: out<=1;
   56056: out<=1;
   56057: out<=1;
   56058: out<=0;
   56059: out<=0;
   56060: out<=1;
   56061: out<=0;
   56062: out<=1;
   56063: out<=0;
   56064: out<=0;
   56065: out<=0;
   56066: out<=1;
   56067: out<=1;
   56068: out<=1;
   56069: out<=0;
   56070: out<=1;
   56071: out<=0;
   56072: out<=0;
   56073: out<=1;
   56074: out<=1;
   56075: out<=0;
   56076: out<=1;
   56077: out<=1;
   56078: out<=1;
   56079: out<=1;
   56080: out<=1;
   56081: out<=0;
   56082: out<=1;
   56083: out<=0;
   56084: out<=1;
   56085: out<=1;
   56086: out<=0;
   56087: out<=0;
   56088: out<=0;
   56089: out<=0;
   56090: out<=0;
   56091: out<=0;
   56092: out<=0;
   56093: out<=1;
   56094: out<=1;
   56095: out<=0;
   56096: out<=1;
   56097: out<=0;
   56098: out<=0;
   56099: out<=1;
   56100: out<=1;
   56101: out<=1;
   56102: out<=1;
   56103: out<=1;
   56104: out<=1;
   56105: out<=1;
   56106: out<=0;
   56107: out<=0;
   56108: out<=1;
   56109: out<=0;
   56110: out<=1;
   56111: out<=0;
   56112: out<=0;
   56113: out<=0;
   56114: out<=0;
   56115: out<=0;
   56116: out<=1;
   56117: out<=0;
   56118: out<=0;
   56119: out<=1;
   56120: out<=1;
   56121: out<=0;
   56122: out<=1;
   56123: out<=0;
   56124: out<=0;
   56125: out<=0;
   56126: out<=1;
   56127: out<=1;
   56128: out<=0;
   56129: out<=0;
   56130: out<=1;
   56131: out<=1;
   56132: out<=1;
   56133: out<=0;
   56134: out<=1;
   56135: out<=0;
   56136: out<=0;
   56137: out<=1;
   56138: out<=1;
   56139: out<=0;
   56140: out<=1;
   56141: out<=1;
   56142: out<=1;
   56143: out<=1;
   56144: out<=0;
   56145: out<=1;
   56146: out<=0;
   56147: out<=1;
   56148: out<=0;
   56149: out<=0;
   56150: out<=1;
   56151: out<=1;
   56152: out<=1;
   56153: out<=1;
   56154: out<=1;
   56155: out<=1;
   56156: out<=1;
   56157: out<=0;
   56158: out<=0;
   56159: out<=1;
   56160: out<=0;
   56161: out<=1;
   56162: out<=1;
   56163: out<=0;
   56164: out<=0;
   56165: out<=0;
   56166: out<=0;
   56167: out<=0;
   56168: out<=0;
   56169: out<=0;
   56170: out<=1;
   56171: out<=1;
   56172: out<=0;
   56173: out<=1;
   56174: out<=0;
   56175: out<=1;
   56176: out<=0;
   56177: out<=0;
   56178: out<=0;
   56179: out<=0;
   56180: out<=1;
   56181: out<=0;
   56182: out<=0;
   56183: out<=1;
   56184: out<=1;
   56185: out<=0;
   56186: out<=1;
   56187: out<=0;
   56188: out<=0;
   56189: out<=0;
   56190: out<=1;
   56191: out<=1;
   56192: out<=0;
   56193: out<=0;
   56194: out<=1;
   56195: out<=1;
   56196: out<=1;
   56197: out<=0;
   56198: out<=1;
   56199: out<=0;
   56200: out<=0;
   56201: out<=1;
   56202: out<=1;
   56203: out<=0;
   56204: out<=1;
   56205: out<=1;
   56206: out<=1;
   56207: out<=1;
   56208: out<=0;
   56209: out<=1;
   56210: out<=0;
   56211: out<=1;
   56212: out<=0;
   56213: out<=0;
   56214: out<=1;
   56215: out<=1;
   56216: out<=1;
   56217: out<=1;
   56218: out<=1;
   56219: out<=1;
   56220: out<=1;
   56221: out<=0;
   56222: out<=0;
   56223: out<=1;
   56224: out<=1;
   56225: out<=0;
   56226: out<=0;
   56227: out<=1;
   56228: out<=1;
   56229: out<=1;
   56230: out<=1;
   56231: out<=1;
   56232: out<=1;
   56233: out<=1;
   56234: out<=0;
   56235: out<=0;
   56236: out<=1;
   56237: out<=0;
   56238: out<=1;
   56239: out<=0;
   56240: out<=1;
   56241: out<=1;
   56242: out<=1;
   56243: out<=1;
   56244: out<=0;
   56245: out<=1;
   56246: out<=1;
   56247: out<=0;
   56248: out<=0;
   56249: out<=1;
   56250: out<=0;
   56251: out<=1;
   56252: out<=1;
   56253: out<=1;
   56254: out<=0;
   56255: out<=0;
   56256: out<=0;
   56257: out<=0;
   56258: out<=1;
   56259: out<=1;
   56260: out<=1;
   56261: out<=0;
   56262: out<=1;
   56263: out<=0;
   56264: out<=0;
   56265: out<=1;
   56266: out<=1;
   56267: out<=0;
   56268: out<=1;
   56269: out<=1;
   56270: out<=1;
   56271: out<=1;
   56272: out<=1;
   56273: out<=0;
   56274: out<=1;
   56275: out<=0;
   56276: out<=1;
   56277: out<=1;
   56278: out<=0;
   56279: out<=0;
   56280: out<=0;
   56281: out<=0;
   56282: out<=0;
   56283: out<=0;
   56284: out<=0;
   56285: out<=1;
   56286: out<=1;
   56287: out<=0;
   56288: out<=0;
   56289: out<=1;
   56290: out<=1;
   56291: out<=0;
   56292: out<=0;
   56293: out<=0;
   56294: out<=0;
   56295: out<=0;
   56296: out<=0;
   56297: out<=0;
   56298: out<=1;
   56299: out<=1;
   56300: out<=0;
   56301: out<=1;
   56302: out<=0;
   56303: out<=1;
   56304: out<=1;
   56305: out<=1;
   56306: out<=1;
   56307: out<=1;
   56308: out<=0;
   56309: out<=1;
   56310: out<=1;
   56311: out<=0;
   56312: out<=0;
   56313: out<=1;
   56314: out<=0;
   56315: out<=1;
   56316: out<=1;
   56317: out<=1;
   56318: out<=0;
   56319: out<=0;
   56320: out<=0;
   56321: out<=1;
   56322: out<=1;
   56323: out<=0;
   56324: out<=1;
   56325: out<=1;
   56326: out<=1;
   56327: out<=1;
   56328: out<=1;
   56329: out<=1;
   56330: out<=0;
   56331: out<=0;
   56332: out<=0;
   56333: out<=1;
   56334: out<=0;
   56335: out<=1;
   56336: out<=1;
   56337: out<=1;
   56338: out<=1;
   56339: out<=1;
   56340: out<=1;
   56341: out<=0;
   56342: out<=0;
   56343: out<=1;
   56344: out<=1;
   56345: out<=0;
   56346: out<=1;
   56347: out<=0;
   56348: out<=1;
   56349: out<=1;
   56350: out<=0;
   56351: out<=0;
   56352: out<=0;
   56353: out<=0;
   56354: out<=1;
   56355: out<=1;
   56356: out<=0;
   56357: out<=1;
   56358: out<=0;
   56359: out<=1;
   56360: out<=1;
   56361: out<=0;
   56362: out<=0;
   56363: out<=1;
   56364: out<=1;
   56365: out<=1;
   56366: out<=1;
   56367: out<=1;
   56368: out<=1;
   56369: out<=0;
   56370: out<=1;
   56371: out<=0;
   56372: out<=0;
   56373: out<=0;
   56374: out<=1;
   56375: out<=1;
   56376: out<=1;
   56377: out<=1;
   56378: out<=1;
   56379: out<=1;
   56380: out<=0;
   56381: out<=1;
   56382: out<=1;
   56383: out<=0;
   56384: out<=1;
   56385: out<=0;
   56386: out<=0;
   56387: out<=1;
   56388: out<=0;
   56389: out<=0;
   56390: out<=0;
   56391: out<=0;
   56392: out<=0;
   56393: out<=0;
   56394: out<=1;
   56395: out<=1;
   56396: out<=1;
   56397: out<=0;
   56398: out<=1;
   56399: out<=0;
   56400: out<=1;
   56401: out<=1;
   56402: out<=1;
   56403: out<=1;
   56404: out<=1;
   56405: out<=0;
   56406: out<=0;
   56407: out<=1;
   56408: out<=1;
   56409: out<=0;
   56410: out<=1;
   56411: out<=0;
   56412: out<=1;
   56413: out<=1;
   56414: out<=0;
   56415: out<=0;
   56416: out<=0;
   56417: out<=0;
   56418: out<=1;
   56419: out<=1;
   56420: out<=0;
   56421: out<=1;
   56422: out<=0;
   56423: out<=1;
   56424: out<=1;
   56425: out<=0;
   56426: out<=0;
   56427: out<=1;
   56428: out<=1;
   56429: out<=1;
   56430: out<=1;
   56431: out<=1;
   56432: out<=0;
   56433: out<=1;
   56434: out<=0;
   56435: out<=1;
   56436: out<=1;
   56437: out<=1;
   56438: out<=0;
   56439: out<=0;
   56440: out<=0;
   56441: out<=0;
   56442: out<=0;
   56443: out<=0;
   56444: out<=1;
   56445: out<=0;
   56446: out<=0;
   56447: out<=1;
   56448: out<=0;
   56449: out<=1;
   56450: out<=1;
   56451: out<=0;
   56452: out<=1;
   56453: out<=1;
   56454: out<=1;
   56455: out<=1;
   56456: out<=1;
   56457: out<=1;
   56458: out<=0;
   56459: out<=0;
   56460: out<=0;
   56461: out<=1;
   56462: out<=0;
   56463: out<=1;
   56464: out<=0;
   56465: out<=0;
   56466: out<=0;
   56467: out<=0;
   56468: out<=0;
   56469: out<=1;
   56470: out<=1;
   56471: out<=0;
   56472: out<=0;
   56473: out<=1;
   56474: out<=0;
   56475: out<=1;
   56476: out<=0;
   56477: out<=0;
   56478: out<=1;
   56479: out<=1;
   56480: out<=0;
   56481: out<=0;
   56482: out<=1;
   56483: out<=1;
   56484: out<=0;
   56485: out<=1;
   56486: out<=0;
   56487: out<=1;
   56488: out<=1;
   56489: out<=0;
   56490: out<=0;
   56491: out<=1;
   56492: out<=1;
   56493: out<=1;
   56494: out<=1;
   56495: out<=1;
   56496: out<=0;
   56497: out<=1;
   56498: out<=0;
   56499: out<=1;
   56500: out<=1;
   56501: out<=1;
   56502: out<=0;
   56503: out<=0;
   56504: out<=0;
   56505: out<=0;
   56506: out<=0;
   56507: out<=0;
   56508: out<=1;
   56509: out<=0;
   56510: out<=0;
   56511: out<=1;
   56512: out<=1;
   56513: out<=0;
   56514: out<=0;
   56515: out<=1;
   56516: out<=0;
   56517: out<=0;
   56518: out<=0;
   56519: out<=0;
   56520: out<=0;
   56521: out<=0;
   56522: out<=1;
   56523: out<=1;
   56524: out<=1;
   56525: out<=0;
   56526: out<=1;
   56527: out<=0;
   56528: out<=0;
   56529: out<=0;
   56530: out<=0;
   56531: out<=0;
   56532: out<=0;
   56533: out<=1;
   56534: out<=1;
   56535: out<=0;
   56536: out<=0;
   56537: out<=1;
   56538: out<=0;
   56539: out<=1;
   56540: out<=0;
   56541: out<=0;
   56542: out<=1;
   56543: out<=1;
   56544: out<=0;
   56545: out<=0;
   56546: out<=1;
   56547: out<=1;
   56548: out<=0;
   56549: out<=1;
   56550: out<=0;
   56551: out<=1;
   56552: out<=1;
   56553: out<=0;
   56554: out<=0;
   56555: out<=1;
   56556: out<=1;
   56557: out<=1;
   56558: out<=1;
   56559: out<=1;
   56560: out<=1;
   56561: out<=0;
   56562: out<=1;
   56563: out<=0;
   56564: out<=0;
   56565: out<=0;
   56566: out<=1;
   56567: out<=1;
   56568: out<=1;
   56569: out<=1;
   56570: out<=1;
   56571: out<=1;
   56572: out<=0;
   56573: out<=1;
   56574: out<=1;
   56575: out<=0;
   56576: out<=1;
   56577: out<=1;
   56578: out<=1;
   56579: out<=1;
   56580: out<=1;
   56581: out<=0;
   56582: out<=0;
   56583: out<=1;
   56584: out<=1;
   56585: out<=0;
   56586: out<=1;
   56587: out<=0;
   56588: out<=1;
   56589: out<=1;
   56590: out<=0;
   56591: out<=0;
   56592: out<=1;
   56593: out<=0;
   56594: out<=0;
   56595: out<=1;
   56596: out<=0;
   56597: out<=0;
   56598: out<=0;
   56599: out<=0;
   56600: out<=0;
   56601: out<=0;
   56602: out<=1;
   56603: out<=1;
   56604: out<=1;
   56605: out<=0;
   56606: out<=1;
   56607: out<=0;
   56608: out<=0;
   56609: out<=1;
   56610: out<=0;
   56611: out<=1;
   56612: out<=1;
   56613: out<=1;
   56614: out<=0;
   56615: out<=0;
   56616: out<=0;
   56617: out<=0;
   56618: out<=0;
   56619: out<=0;
   56620: out<=1;
   56621: out<=0;
   56622: out<=0;
   56623: out<=1;
   56624: out<=0;
   56625: out<=0;
   56626: out<=1;
   56627: out<=1;
   56628: out<=0;
   56629: out<=1;
   56630: out<=0;
   56631: out<=1;
   56632: out<=1;
   56633: out<=0;
   56634: out<=0;
   56635: out<=1;
   56636: out<=1;
   56637: out<=1;
   56638: out<=1;
   56639: out<=1;
   56640: out<=1;
   56641: out<=1;
   56642: out<=1;
   56643: out<=1;
   56644: out<=1;
   56645: out<=0;
   56646: out<=0;
   56647: out<=1;
   56648: out<=1;
   56649: out<=0;
   56650: out<=1;
   56651: out<=0;
   56652: out<=1;
   56653: out<=1;
   56654: out<=0;
   56655: out<=0;
   56656: out<=0;
   56657: out<=1;
   56658: out<=1;
   56659: out<=0;
   56660: out<=1;
   56661: out<=1;
   56662: out<=1;
   56663: out<=1;
   56664: out<=1;
   56665: out<=1;
   56666: out<=0;
   56667: out<=0;
   56668: out<=0;
   56669: out<=1;
   56670: out<=0;
   56671: out<=1;
   56672: out<=1;
   56673: out<=0;
   56674: out<=1;
   56675: out<=0;
   56676: out<=0;
   56677: out<=0;
   56678: out<=1;
   56679: out<=1;
   56680: out<=1;
   56681: out<=1;
   56682: out<=1;
   56683: out<=1;
   56684: out<=0;
   56685: out<=1;
   56686: out<=1;
   56687: out<=0;
   56688: out<=0;
   56689: out<=0;
   56690: out<=1;
   56691: out<=1;
   56692: out<=0;
   56693: out<=1;
   56694: out<=0;
   56695: out<=1;
   56696: out<=1;
   56697: out<=0;
   56698: out<=0;
   56699: out<=1;
   56700: out<=1;
   56701: out<=1;
   56702: out<=1;
   56703: out<=1;
   56704: out<=0;
   56705: out<=0;
   56706: out<=0;
   56707: out<=0;
   56708: out<=0;
   56709: out<=1;
   56710: out<=1;
   56711: out<=0;
   56712: out<=0;
   56713: out<=1;
   56714: out<=0;
   56715: out<=1;
   56716: out<=0;
   56717: out<=0;
   56718: out<=1;
   56719: out<=1;
   56720: out<=1;
   56721: out<=0;
   56722: out<=0;
   56723: out<=1;
   56724: out<=0;
   56725: out<=0;
   56726: out<=0;
   56727: out<=0;
   56728: out<=0;
   56729: out<=0;
   56730: out<=1;
   56731: out<=1;
   56732: out<=1;
   56733: out<=0;
   56734: out<=1;
   56735: out<=0;
   56736: out<=1;
   56737: out<=0;
   56738: out<=1;
   56739: out<=0;
   56740: out<=0;
   56741: out<=0;
   56742: out<=1;
   56743: out<=1;
   56744: out<=1;
   56745: out<=1;
   56746: out<=1;
   56747: out<=1;
   56748: out<=0;
   56749: out<=1;
   56750: out<=1;
   56751: out<=0;
   56752: out<=0;
   56753: out<=0;
   56754: out<=1;
   56755: out<=1;
   56756: out<=0;
   56757: out<=1;
   56758: out<=0;
   56759: out<=1;
   56760: out<=1;
   56761: out<=0;
   56762: out<=0;
   56763: out<=1;
   56764: out<=1;
   56765: out<=1;
   56766: out<=1;
   56767: out<=1;
   56768: out<=0;
   56769: out<=0;
   56770: out<=0;
   56771: out<=0;
   56772: out<=0;
   56773: out<=1;
   56774: out<=1;
   56775: out<=0;
   56776: out<=0;
   56777: out<=1;
   56778: out<=0;
   56779: out<=1;
   56780: out<=0;
   56781: out<=0;
   56782: out<=1;
   56783: out<=1;
   56784: out<=0;
   56785: out<=1;
   56786: out<=1;
   56787: out<=0;
   56788: out<=1;
   56789: out<=1;
   56790: out<=1;
   56791: out<=1;
   56792: out<=1;
   56793: out<=1;
   56794: out<=0;
   56795: out<=0;
   56796: out<=0;
   56797: out<=1;
   56798: out<=0;
   56799: out<=1;
   56800: out<=0;
   56801: out<=1;
   56802: out<=0;
   56803: out<=1;
   56804: out<=1;
   56805: out<=1;
   56806: out<=0;
   56807: out<=0;
   56808: out<=0;
   56809: out<=0;
   56810: out<=0;
   56811: out<=0;
   56812: out<=1;
   56813: out<=0;
   56814: out<=0;
   56815: out<=1;
   56816: out<=0;
   56817: out<=0;
   56818: out<=1;
   56819: out<=1;
   56820: out<=0;
   56821: out<=1;
   56822: out<=0;
   56823: out<=1;
   56824: out<=1;
   56825: out<=0;
   56826: out<=0;
   56827: out<=1;
   56828: out<=1;
   56829: out<=1;
   56830: out<=1;
   56831: out<=1;
   56832: out<=0;
   56833: out<=0;
   56834: out<=1;
   56835: out<=1;
   56836: out<=0;
   56837: out<=1;
   56838: out<=0;
   56839: out<=1;
   56840: out<=1;
   56841: out<=0;
   56842: out<=0;
   56843: out<=1;
   56844: out<=1;
   56845: out<=1;
   56846: out<=1;
   56847: out<=1;
   56848: out<=0;
   56849: out<=1;
   56850: out<=0;
   56851: out<=1;
   56852: out<=1;
   56853: out<=1;
   56854: out<=0;
   56855: out<=0;
   56856: out<=0;
   56857: out<=0;
   56858: out<=0;
   56859: out<=0;
   56860: out<=1;
   56861: out<=0;
   56862: out<=0;
   56863: out<=1;
   56864: out<=0;
   56865: out<=1;
   56866: out<=1;
   56867: out<=0;
   56868: out<=1;
   56869: out<=1;
   56870: out<=1;
   56871: out<=1;
   56872: out<=1;
   56873: out<=1;
   56874: out<=0;
   56875: out<=0;
   56876: out<=0;
   56877: out<=1;
   56878: out<=0;
   56879: out<=1;
   56880: out<=0;
   56881: out<=0;
   56882: out<=0;
   56883: out<=0;
   56884: out<=0;
   56885: out<=1;
   56886: out<=1;
   56887: out<=0;
   56888: out<=0;
   56889: out<=1;
   56890: out<=0;
   56891: out<=1;
   56892: out<=0;
   56893: out<=0;
   56894: out<=1;
   56895: out<=1;
   56896: out<=0;
   56897: out<=0;
   56898: out<=1;
   56899: out<=1;
   56900: out<=0;
   56901: out<=1;
   56902: out<=0;
   56903: out<=1;
   56904: out<=1;
   56905: out<=0;
   56906: out<=0;
   56907: out<=1;
   56908: out<=1;
   56909: out<=1;
   56910: out<=1;
   56911: out<=1;
   56912: out<=1;
   56913: out<=0;
   56914: out<=1;
   56915: out<=0;
   56916: out<=0;
   56917: out<=0;
   56918: out<=1;
   56919: out<=1;
   56920: out<=1;
   56921: out<=1;
   56922: out<=1;
   56923: out<=1;
   56924: out<=0;
   56925: out<=1;
   56926: out<=1;
   56927: out<=0;
   56928: out<=1;
   56929: out<=0;
   56930: out<=0;
   56931: out<=1;
   56932: out<=0;
   56933: out<=0;
   56934: out<=0;
   56935: out<=0;
   56936: out<=0;
   56937: out<=0;
   56938: out<=1;
   56939: out<=1;
   56940: out<=1;
   56941: out<=0;
   56942: out<=1;
   56943: out<=0;
   56944: out<=0;
   56945: out<=0;
   56946: out<=0;
   56947: out<=0;
   56948: out<=0;
   56949: out<=1;
   56950: out<=1;
   56951: out<=0;
   56952: out<=0;
   56953: out<=1;
   56954: out<=0;
   56955: out<=1;
   56956: out<=0;
   56957: out<=0;
   56958: out<=1;
   56959: out<=1;
   56960: out<=0;
   56961: out<=0;
   56962: out<=1;
   56963: out<=1;
   56964: out<=0;
   56965: out<=1;
   56966: out<=0;
   56967: out<=1;
   56968: out<=1;
   56969: out<=0;
   56970: out<=0;
   56971: out<=1;
   56972: out<=1;
   56973: out<=1;
   56974: out<=1;
   56975: out<=1;
   56976: out<=1;
   56977: out<=0;
   56978: out<=1;
   56979: out<=0;
   56980: out<=0;
   56981: out<=0;
   56982: out<=1;
   56983: out<=1;
   56984: out<=1;
   56985: out<=1;
   56986: out<=1;
   56987: out<=1;
   56988: out<=0;
   56989: out<=1;
   56990: out<=1;
   56991: out<=0;
   56992: out<=0;
   56993: out<=1;
   56994: out<=1;
   56995: out<=0;
   56996: out<=1;
   56997: out<=1;
   56998: out<=1;
   56999: out<=1;
   57000: out<=1;
   57001: out<=1;
   57002: out<=0;
   57003: out<=0;
   57004: out<=0;
   57005: out<=1;
   57006: out<=0;
   57007: out<=1;
   57008: out<=1;
   57009: out<=1;
   57010: out<=1;
   57011: out<=1;
   57012: out<=1;
   57013: out<=0;
   57014: out<=0;
   57015: out<=1;
   57016: out<=1;
   57017: out<=0;
   57018: out<=1;
   57019: out<=0;
   57020: out<=1;
   57021: out<=1;
   57022: out<=0;
   57023: out<=0;
   57024: out<=0;
   57025: out<=0;
   57026: out<=1;
   57027: out<=1;
   57028: out<=0;
   57029: out<=1;
   57030: out<=0;
   57031: out<=1;
   57032: out<=1;
   57033: out<=0;
   57034: out<=0;
   57035: out<=1;
   57036: out<=1;
   57037: out<=1;
   57038: out<=1;
   57039: out<=1;
   57040: out<=0;
   57041: out<=1;
   57042: out<=0;
   57043: out<=1;
   57044: out<=1;
   57045: out<=1;
   57046: out<=0;
   57047: out<=0;
   57048: out<=0;
   57049: out<=0;
   57050: out<=0;
   57051: out<=0;
   57052: out<=1;
   57053: out<=0;
   57054: out<=0;
   57055: out<=1;
   57056: out<=1;
   57057: out<=0;
   57058: out<=0;
   57059: out<=1;
   57060: out<=0;
   57061: out<=0;
   57062: out<=0;
   57063: out<=0;
   57064: out<=0;
   57065: out<=0;
   57066: out<=1;
   57067: out<=1;
   57068: out<=1;
   57069: out<=0;
   57070: out<=1;
   57071: out<=0;
   57072: out<=1;
   57073: out<=1;
   57074: out<=1;
   57075: out<=1;
   57076: out<=1;
   57077: out<=0;
   57078: out<=0;
   57079: out<=1;
   57080: out<=1;
   57081: out<=0;
   57082: out<=1;
   57083: out<=0;
   57084: out<=1;
   57085: out<=1;
   57086: out<=0;
   57087: out<=0;
   57088: out<=1;
   57089: out<=0;
   57090: out<=1;
   57091: out<=0;
   57092: out<=0;
   57093: out<=0;
   57094: out<=1;
   57095: out<=1;
   57096: out<=1;
   57097: out<=1;
   57098: out<=1;
   57099: out<=1;
   57100: out<=0;
   57101: out<=1;
   57102: out<=1;
   57103: out<=0;
   57104: out<=0;
   57105: out<=0;
   57106: out<=1;
   57107: out<=1;
   57108: out<=0;
   57109: out<=1;
   57110: out<=0;
   57111: out<=1;
   57112: out<=1;
   57113: out<=0;
   57114: out<=0;
   57115: out<=1;
   57116: out<=1;
   57117: out<=1;
   57118: out<=1;
   57119: out<=1;
   57120: out<=0;
   57121: out<=0;
   57122: out<=0;
   57123: out<=0;
   57124: out<=0;
   57125: out<=1;
   57126: out<=1;
   57127: out<=0;
   57128: out<=0;
   57129: out<=1;
   57130: out<=0;
   57131: out<=1;
   57132: out<=0;
   57133: out<=0;
   57134: out<=1;
   57135: out<=1;
   57136: out<=1;
   57137: out<=0;
   57138: out<=0;
   57139: out<=1;
   57140: out<=0;
   57141: out<=0;
   57142: out<=0;
   57143: out<=0;
   57144: out<=0;
   57145: out<=0;
   57146: out<=1;
   57147: out<=1;
   57148: out<=1;
   57149: out<=0;
   57150: out<=1;
   57151: out<=0;
   57152: out<=0;
   57153: out<=1;
   57154: out<=0;
   57155: out<=1;
   57156: out<=1;
   57157: out<=1;
   57158: out<=0;
   57159: out<=0;
   57160: out<=0;
   57161: out<=0;
   57162: out<=0;
   57163: out<=0;
   57164: out<=1;
   57165: out<=0;
   57166: out<=0;
   57167: out<=1;
   57168: out<=0;
   57169: out<=0;
   57170: out<=1;
   57171: out<=1;
   57172: out<=0;
   57173: out<=1;
   57174: out<=0;
   57175: out<=1;
   57176: out<=1;
   57177: out<=0;
   57178: out<=0;
   57179: out<=1;
   57180: out<=1;
   57181: out<=1;
   57182: out<=1;
   57183: out<=1;
   57184: out<=0;
   57185: out<=0;
   57186: out<=0;
   57187: out<=0;
   57188: out<=0;
   57189: out<=1;
   57190: out<=1;
   57191: out<=0;
   57192: out<=0;
   57193: out<=1;
   57194: out<=0;
   57195: out<=1;
   57196: out<=0;
   57197: out<=0;
   57198: out<=1;
   57199: out<=1;
   57200: out<=0;
   57201: out<=1;
   57202: out<=1;
   57203: out<=0;
   57204: out<=1;
   57205: out<=1;
   57206: out<=1;
   57207: out<=1;
   57208: out<=1;
   57209: out<=1;
   57210: out<=0;
   57211: out<=0;
   57212: out<=0;
   57213: out<=1;
   57214: out<=0;
   57215: out<=1;
   57216: out<=0;
   57217: out<=1;
   57218: out<=0;
   57219: out<=1;
   57220: out<=1;
   57221: out<=1;
   57222: out<=0;
   57223: out<=0;
   57224: out<=0;
   57225: out<=0;
   57226: out<=0;
   57227: out<=0;
   57228: out<=1;
   57229: out<=0;
   57230: out<=0;
   57231: out<=1;
   57232: out<=0;
   57233: out<=0;
   57234: out<=1;
   57235: out<=1;
   57236: out<=0;
   57237: out<=1;
   57238: out<=0;
   57239: out<=1;
   57240: out<=1;
   57241: out<=0;
   57242: out<=0;
   57243: out<=1;
   57244: out<=1;
   57245: out<=1;
   57246: out<=1;
   57247: out<=1;
   57248: out<=1;
   57249: out<=1;
   57250: out<=1;
   57251: out<=1;
   57252: out<=1;
   57253: out<=0;
   57254: out<=0;
   57255: out<=1;
   57256: out<=1;
   57257: out<=0;
   57258: out<=1;
   57259: out<=0;
   57260: out<=1;
   57261: out<=1;
   57262: out<=0;
   57263: out<=0;
   57264: out<=1;
   57265: out<=0;
   57266: out<=0;
   57267: out<=1;
   57268: out<=0;
   57269: out<=0;
   57270: out<=0;
   57271: out<=0;
   57272: out<=0;
   57273: out<=0;
   57274: out<=1;
   57275: out<=1;
   57276: out<=1;
   57277: out<=0;
   57278: out<=1;
   57279: out<=0;
   57280: out<=1;
   57281: out<=0;
   57282: out<=1;
   57283: out<=0;
   57284: out<=0;
   57285: out<=0;
   57286: out<=1;
   57287: out<=1;
   57288: out<=1;
   57289: out<=1;
   57290: out<=1;
   57291: out<=1;
   57292: out<=0;
   57293: out<=1;
   57294: out<=1;
   57295: out<=0;
   57296: out<=0;
   57297: out<=0;
   57298: out<=1;
   57299: out<=1;
   57300: out<=0;
   57301: out<=1;
   57302: out<=0;
   57303: out<=1;
   57304: out<=1;
   57305: out<=0;
   57306: out<=0;
   57307: out<=1;
   57308: out<=1;
   57309: out<=1;
   57310: out<=1;
   57311: out<=1;
   57312: out<=1;
   57313: out<=1;
   57314: out<=1;
   57315: out<=1;
   57316: out<=1;
   57317: out<=0;
   57318: out<=0;
   57319: out<=1;
   57320: out<=1;
   57321: out<=0;
   57322: out<=1;
   57323: out<=0;
   57324: out<=1;
   57325: out<=1;
   57326: out<=0;
   57327: out<=0;
   57328: out<=0;
   57329: out<=1;
   57330: out<=1;
   57331: out<=0;
   57332: out<=1;
   57333: out<=1;
   57334: out<=1;
   57335: out<=1;
   57336: out<=1;
   57337: out<=1;
   57338: out<=0;
   57339: out<=0;
   57340: out<=0;
   57341: out<=1;
   57342: out<=0;
   57343: out<=1;
   57344: out<=0;
   57345: out<=1;
   57346: out<=0;
   57347: out<=1;
   57348: out<=1;
   57349: out<=1;
   57350: out<=0;
   57351: out<=0;
   57352: out<=0;
   57353: out<=0;
   57354: out<=0;
   57355: out<=0;
   57356: out<=1;
   57357: out<=0;
   57358: out<=0;
   57359: out<=1;
   57360: out<=1;
   57361: out<=1;
   57362: out<=0;
   57363: out<=0;
   57364: out<=1;
   57365: out<=0;
   57366: out<=1;
   57367: out<=0;
   57368: out<=0;
   57369: out<=1;
   57370: out<=1;
   57371: out<=0;
   57372: out<=0;
   57373: out<=0;
   57374: out<=0;
   57375: out<=0;
   57376: out<=0;
   57377: out<=0;
   57378: out<=0;
   57379: out<=0;
   57380: out<=0;
   57381: out<=1;
   57382: out<=1;
   57383: out<=0;
   57384: out<=0;
   57385: out<=1;
   57386: out<=0;
   57387: out<=1;
   57388: out<=0;
   57389: out<=0;
   57390: out<=1;
   57391: out<=1;
   57392: out<=1;
   57393: out<=0;
   57394: out<=0;
   57395: out<=1;
   57396: out<=0;
   57397: out<=0;
   57398: out<=0;
   57399: out<=0;
   57400: out<=0;
   57401: out<=0;
   57402: out<=1;
   57403: out<=1;
   57404: out<=1;
   57405: out<=0;
   57406: out<=1;
   57407: out<=0;
   57408: out<=1;
   57409: out<=0;
   57410: out<=1;
   57411: out<=0;
   57412: out<=0;
   57413: out<=0;
   57414: out<=1;
   57415: out<=1;
   57416: out<=1;
   57417: out<=1;
   57418: out<=1;
   57419: out<=1;
   57420: out<=0;
   57421: out<=1;
   57422: out<=1;
   57423: out<=0;
   57424: out<=1;
   57425: out<=1;
   57426: out<=0;
   57427: out<=0;
   57428: out<=1;
   57429: out<=0;
   57430: out<=1;
   57431: out<=0;
   57432: out<=0;
   57433: out<=1;
   57434: out<=1;
   57435: out<=0;
   57436: out<=0;
   57437: out<=0;
   57438: out<=0;
   57439: out<=0;
   57440: out<=0;
   57441: out<=0;
   57442: out<=0;
   57443: out<=0;
   57444: out<=0;
   57445: out<=1;
   57446: out<=1;
   57447: out<=0;
   57448: out<=0;
   57449: out<=1;
   57450: out<=0;
   57451: out<=1;
   57452: out<=0;
   57453: out<=0;
   57454: out<=1;
   57455: out<=1;
   57456: out<=0;
   57457: out<=1;
   57458: out<=1;
   57459: out<=0;
   57460: out<=1;
   57461: out<=1;
   57462: out<=1;
   57463: out<=1;
   57464: out<=1;
   57465: out<=1;
   57466: out<=0;
   57467: out<=0;
   57468: out<=0;
   57469: out<=1;
   57470: out<=0;
   57471: out<=1;
   57472: out<=1;
   57473: out<=0;
   57474: out<=1;
   57475: out<=0;
   57476: out<=0;
   57477: out<=0;
   57478: out<=1;
   57479: out<=1;
   57480: out<=1;
   57481: out<=1;
   57482: out<=1;
   57483: out<=1;
   57484: out<=0;
   57485: out<=1;
   57486: out<=1;
   57487: out<=0;
   57488: out<=1;
   57489: out<=1;
   57490: out<=0;
   57491: out<=0;
   57492: out<=1;
   57493: out<=0;
   57494: out<=1;
   57495: out<=0;
   57496: out<=0;
   57497: out<=1;
   57498: out<=1;
   57499: out<=0;
   57500: out<=0;
   57501: out<=0;
   57502: out<=0;
   57503: out<=0;
   57504: out<=1;
   57505: out<=1;
   57506: out<=1;
   57507: out<=1;
   57508: out<=1;
   57509: out<=0;
   57510: out<=0;
   57511: out<=1;
   57512: out<=1;
   57513: out<=0;
   57514: out<=1;
   57515: out<=0;
   57516: out<=1;
   57517: out<=1;
   57518: out<=0;
   57519: out<=0;
   57520: out<=1;
   57521: out<=0;
   57522: out<=0;
   57523: out<=1;
   57524: out<=0;
   57525: out<=0;
   57526: out<=0;
   57527: out<=0;
   57528: out<=0;
   57529: out<=0;
   57530: out<=1;
   57531: out<=1;
   57532: out<=1;
   57533: out<=0;
   57534: out<=1;
   57535: out<=0;
   57536: out<=0;
   57537: out<=1;
   57538: out<=0;
   57539: out<=1;
   57540: out<=1;
   57541: out<=1;
   57542: out<=0;
   57543: out<=0;
   57544: out<=0;
   57545: out<=0;
   57546: out<=0;
   57547: out<=0;
   57548: out<=1;
   57549: out<=0;
   57550: out<=0;
   57551: out<=1;
   57552: out<=1;
   57553: out<=1;
   57554: out<=0;
   57555: out<=0;
   57556: out<=1;
   57557: out<=0;
   57558: out<=1;
   57559: out<=0;
   57560: out<=0;
   57561: out<=1;
   57562: out<=1;
   57563: out<=0;
   57564: out<=0;
   57565: out<=0;
   57566: out<=0;
   57567: out<=0;
   57568: out<=1;
   57569: out<=1;
   57570: out<=1;
   57571: out<=1;
   57572: out<=1;
   57573: out<=0;
   57574: out<=0;
   57575: out<=1;
   57576: out<=1;
   57577: out<=0;
   57578: out<=1;
   57579: out<=0;
   57580: out<=1;
   57581: out<=1;
   57582: out<=0;
   57583: out<=0;
   57584: out<=0;
   57585: out<=1;
   57586: out<=1;
   57587: out<=0;
   57588: out<=1;
   57589: out<=1;
   57590: out<=1;
   57591: out<=1;
   57592: out<=1;
   57593: out<=1;
   57594: out<=0;
   57595: out<=0;
   57596: out<=0;
   57597: out<=1;
   57598: out<=0;
   57599: out<=1;
   57600: out<=1;
   57601: out<=1;
   57602: out<=0;
   57603: out<=0;
   57604: out<=1;
   57605: out<=0;
   57606: out<=1;
   57607: out<=0;
   57608: out<=0;
   57609: out<=1;
   57610: out<=1;
   57611: out<=0;
   57612: out<=0;
   57613: out<=0;
   57614: out<=0;
   57615: out<=0;
   57616: out<=1;
   57617: out<=0;
   57618: out<=1;
   57619: out<=0;
   57620: out<=0;
   57621: out<=0;
   57622: out<=1;
   57623: out<=1;
   57624: out<=1;
   57625: out<=1;
   57626: out<=1;
   57627: out<=1;
   57628: out<=0;
   57629: out<=1;
   57630: out<=1;
   57631: out<=0;
   57632: out<=0;
   57633: out<=1;
   57634: out<=1;
   57635: out<=0;
   57636: out<=1;
   57637: out<=1;
   57638: out<=1;
   57639: out<=1;
   57640: out<=1;
   57641: out<=1;
   57642: out<=0;
   57643: out<=0;
   57644: out<=0;
   57645: out<=1;
   57646: out<=0;
   57647: out<=1;
   57648: out<=0;
   57649: out<=0;
   57650: out<=0;
   57651: out<=0;
   57652: out<=0;
   57653: out<=1;
   57654: out<=1;
   57655: out<=0;
   57656: out<=0;
   57657: out<=1;
   57658: out<=0;
   57659: out<=1;
   57660: out<=0;
   57661: out<=0;
   57662: out<=1;
   57663: out<=1;
   57664: out<=1;
   57665: out<=1;
   57666: out<=0;
   57667: out<=0;
   57668: out<=1;
   57669: out<=0;
   57670: out<=1;
   57671: out<=0;
   57672: out<=0;
   57673: out<=1;
   57674: out<=1;
   57675: out<=0;
   57676: out<=0;
   57677: out<=0;
   57678: out<=0;
   57679: out<=0;
   57680: out<=0;
   57681: out<=1;
   57682: out<=0;
   57683: out<=1;
   57684: out<=1;
   57685: out<=1;
   57686: out<=0;
   57687: out<=0;
   57688: out<=0;
   57689: out<=0;
   57690: out<=0;
   57691: out<=0;
   57692: out<=1;
   57693: out<=0;
   57694: out<=0;
   57695: out<=1;
   57696: out<=1;
   57697: out<=0;
   57698: out<=0;
   57699: out<=1;
   57700: out<=0;
   57701: out<=0;
   57702: out<=0;
   57703: out<=0;
   57704: out<=0;
   57705: out<=0;
   57706: out<=1;
   57707: out<=1;
   57708: out<=1;
   57709: out<=0;
   57710: out<=1;
   57711: out<=0;
   57712: out<=0;
   57713: out<=0;
   57714: out<=0;
   57715: out<=0;
   57716: out<=0;
   57717: out<=1;
   57718: out<=1;
   57719: out<=0;
   57720: out<=0;
   57721: out<=1;
   57722: out<=0;
   57723: out<=1;
   57724: out<=0;
   57725: out<=0;
   57726: out<=1;
   57727: out<=1;
   57728: out<=1;
   57729: out<=1;
   57730: out<=0;
   57731: out<=0;
   57732: out<=1;
   57733: out<=0;
   57734: out<=1;
   57735: out<=0;
   57736: out<=0;
   57737: out<=1;
   57738: out<=1;
   57739: out<=0;
   57740: out<=0;
   57741: out<=0;
   57742: out<=0;
   57743: out<=0;
   57744: out<=0;
   57745: out<=1;
   57746: out<=0;
   57747: out<=1;
   57748: out<=1;
   57749: out<=1;
   57750: out<=0;
   57751: out<=0;
   57752: out<=0;
   57753: out<=0;
   57754: out<=0;
   57755: out<=0;
   57756: out<=1;
   57757: out<=0;
   57758: out<=0;
   57759: out<=1;
   57760: out<=0;
   57761: out<=1;
   57762: out<=1;
   57763: out<=0;
   57764: out<=1;
   57765: out<=1;
   57766: out<=1;
   57767: out<=1;
   57768: out<=1;
   57769: out<=1;
   57770: out<=0;
   57771: out<=0;
   57772: out<=0;
   57773: out<=1;
   57774: out<=0;
   57775: out<=1;
   57776: out<=1;
   57777: out<=1;
   57778: out<=1;
   57779: out<=1;
   57780: out<=1;
   57781: out<=0;
   57782: out<=0;
   57783: out<=1;
   57784: out<=1;
   57785: out<=0;
   57786: out<=1;
   57787: out<=0;
   57788: out<=1;
   57789: out<=1;
   57790: out<=0;
   57791: out<=0;
   57792: out<=1;
   57793: out<=1;
   57794: out<=0;
   57795: out<=0;
   57796: out<=1;
   57797: out<=0;
   57798: out<=1;
   57799: out<=0;
   57800: out<=0;
   57801: out<=1;
   57802: out<=1;
   57803: out<=0;
   57804: out<=0;
   57805: out<=0;
   57806: out<=0;
   57807: out<=0;
   57808: out<=1;
   57809: out<=0;
   57810: out<=1;
   57811: out<=0;
   57812: out<=0;
   57813: out<=0;
   57814: out<=1;
   57815: out<=1;
   57816: out<=1;
   57817: out<=1;
   57818: out<=1;
   57819: out<=1;
   57820: out<=0;
   57821: out<=1;
   57822: out<=1;
   57823: out<=0;
   57824: out<=1;
   57825: out<=0;
   57826: out<=0;
   57827: out<=1;
   57828: out<=0;
   57829: out<=0;
   57830: out<=0;
   57831: out<=0;
   57832: out<=0;
   57833: out<=0;
   57834: out<=1;
   57835: out<=1;
   57836: out<=1;
   57837: out<=0;
   57838: out<=1;
   57839: out<=0;
   57840: out<=1;
   57841: out<=1;
   57842: out<=1;
   57843: out<=1;
   57844: out<=1;
   57845: out<=0;
   57846: out<=0;
   57847: out<=1;
   57848: out<=1;
   57849: out<=0;
   57850: out<=1;
   57851: out<=0;
   57852: out<=1;
   57853: out<=1;
   57854: out<=0;
   57855: out<=0;
   57856: out<=1;
   57857: out<=1;
   57858: out<=1;
   57859: out<=1;
   57860: out<=1;
   57861: out<=0;
   57862: out<=0;
   57863: out<=1;
   57864: out<=1;
   57865: out<=0;
   57866: out<=1;
   57867: out<=0;
   57868: out<=1;
   57869: out<=1;
   57870: out<=0;
   57871: out<=0;
   57872: out<=1;
   57873: out<=0;
   57874: out<=0;
   57875: out<=1;
   57876: out<=0;
   57877: out<=0;
   57878: out<=0;
   57879: out<=0;
   57880: out<=0;
   57881: out<=0;
   57882: out<=1;
   57883: out<=1;
   57884: out<=1;
   57885: out<=0;
   57886: out<=1;
   57887: out<=0;
   57888: out<=1;
   57889: out<=0;
   57890: out<=1;
   57891: out<=0;
   57892: out<=0;
   57893: out<=0;
   57894: out<=1;
   57895: out<=1;
   57896: out<=1;
   57897: out<=1;
   57898: out<=1;
   57899: out<=1;
   57900: out<=0;
   57901: out<=1;
   57902: out<=1;
   57903: out<=0;
   57904: out<=1;
   57905: out<=1;
   57906: out<=0;
   57907: out<=0;
   57908: out<=1;
   57909: out<=0;
   57910: out<=1;
   57911: out<=0;
   57912: out<=0;
   57913: out<=1;
   57914: out<=1;
   57915: out<=0;
   57916: out<=0;
   57917: out<=0;
   57918: out<=0;
   57919: out<=0;
   57920: out<=1;
   57921: out<=1;
   57922: out<=1;
   57923: out<=1;
   57924: out<=1;
   57925: out<=0;
   57926: out<=0;
   57927: out<=1;
   57928: out<=1;
   57929: out<=0;
   57930: out<=1;
   57931: out<=0;
   57932: out<=1;
   57933: out<=1;
   57934: out<=0;
   57935: out<=0;
   57936: out<=0;
   57937: out<=1;
   57938: out<=1;
   57939: out<=0;
   57940: out<=1;
   57941: out<=1;
   57942: out<=1;
   57943: out<=1;
   57944: out<=1;
   57945: out<=1;
   57946: out<=0;
   57947: out<=0;
   57948: out<=0;
   57949: out<=1;
   57950: out<=0;
   57951: out<=1;
   57952: out<=0;
   57953: out<=1;
   57954: out<=0;
   57955: out<=1;
   57956: out<=1;
   57957: out<=1;
   57958: out<=0;
   57959: out<=0;
   57960: out<=0;
   57961: out<=0;
   57962: out<=0;
   57963: out<=0;
   57964: out<=1;
   57965: out<=0;
   57966: out<=0;
   57967: out<=1;
   57968: out<=1;
   57969: out<=1;
   57970: out<=0;
   57971: out<=0;
   57972: out<=1;
   57973: out<=0;
   57974: out<=1;
   57975: out<=0;
   57976: out<=0;
   57977: out<=1;
   57978: out<=1;
   57979: out<=0;
   57980: out<=0;
   57981: out<=0;
   57982: out<=0;
   57983: out<=0;
   57984: out<=0;
   57985: out<=0;
   57986: out<=0;
   57987: out<=0;
   57988: out<=0;
   57989: out<=1;
   57990: out<=1;
   57991: out<=0;
   57992: out<=0;
   57993: out<=1;
   57994: out<=0;
   57995: out<=1;
   57996: out<=0;
   57997: out<=0;
   57998: out<=1;
   57999: out<=1;
   58000: out<=1;
   58001: out<=0;
   58002: out<=0;
   58003: out<=1;
   58004: out<=0;
   58005: out<=0;
   58006: out<=0;
   58007: out<=0;
   58008: out<=0;
   58009: out<=0;
   58010: out<=1;
   58011: out<=1;
   58012: out<=1;
   58013: out<=0;
   58014: out<=1;
   58015: out<=0;
   58016: out<=0;
   58017: out<=1;
   58018: out<=0;
   58019: out<=1;
   58020: out<=1;
   58021: out<=1;
   58022: out<=0;
   58023: out<=0;
   58024: out<=0;
   58025: out<=0;
   58026: out<=0;
   58027: out<=0;
   58028: out<=1;
   58029: out<=0;
   58030: out<=0;
   58031: out<=1;
   58032: out<=1;
   58033: out<=1;
   58034: out<=0;
   58035: out<=0;
   58036: out<=1;
   58037: out<=0;
   58038: out<=1;
   58039: out<=0;
   58040: out<=0;
   58041: out<=1;
   58042: out<=1;
   58043: out<=0;
   58044: out<=0;
   58045: out<=0;
   58046: out<=0;
   58047: out<=0;
   58048: out<=0;
   58049: out<=0;
   58050: out<=0;
   58051: out<=0;
   58052: out<=0;
   58053: out<=1;
   58054: out<=1;
   58055: out<=0;
   58056: out<=0;
   58057: out<=1;
   58058: out<=0;
   58059: out<=1;
   58060: out<=0;
   58061: out<=0;
   58062: out<=1;
   58063: out<=1;
   58064: out<=0;
   58065: out<=1;
   58066: out<=1;
   58067: out<=0;
   58068: out<=1;
   58069: out<=1;
   58070: out<=1;
   58071: out<=1;
   58072: out<=1;
   58073: out<=1;
   58074: out<=0;
   58075: out<=0;
   58076: out<=0;
   58077: out<=1;
   58078: out<=0;
   58079: out<=1;
   58080: out<=1;
   58081: out<=0;
   58082: out<=1;
   58083: out<=0;
   58084: out<=0;
   58085: out<=0;
   58086: out<=1;
   58087: out<=1;
   58088: out<=1;
   58089: out<=1;
   58090: out<=1;
   58091: out<=1;
   58092: out<=0;
   58093: out<=1;
   58094: out<=1;
   58095: out<=0;
   58096: out<=1;
   58097: out<=1;
   58098: out<=0;
   58099: out<=0;
   58100: out<=1;
   58101: out<=0;
   58102: out<=1;
   58103: out<=0;
   58104: out<=0;
   58105: out<=1;
   58106: out<=1;
   58107: out<=0;
   58108: out<=0;
   58109: out<=0;
   58110: out<=0;
   58111: out<=0;
   58112: out<=0;
   58113: out<=1;
   58114: out<=1;
   58115: out<=0;
   58116: out<=1;
   58117: out<=1;
   58118: out<=1;
   58119: out<=1;
   58120: out<=1;
   58121: out<=1;
   58122: out<=0;
   58123: out<=0;
   58124: out<=0;
   58125: out<=1;
   58126: out<=0;
   58127: out<=1;
   58128: out<=1;
   58129: out<=1;
   58130: out<=1;
   58131: out<=1;
   58132: out<=1;
   58133: out<=0;
   58134: out<=0;
   58135: out<=1;
   58136: out<=1;
   58137: out<=0;
   58138: out<=1;
   58139: out<=0;
   58140: out<=1;
   58141: out<=1;
   58142: out<=0;
   58143: out<=0;
   58144: out<=1;
   58145: out<=1;
   58146: out<=0;
   58147: out<=0;
   58148: out<=1;
   58149: out<=0;
   58150: out<=1;
   58151: out<=0;
   58152: out<=0;
   58153: out<=1;
   58154: out<=1;
   58155: out<=0;
   58156: out<=0;
   58157: out<=0;
   58158: out<=0;
   58159: out<=0;
   58160: out<=0;
   58161: out<=1;
   58162: out<=0;
   58163: out<=1;
   58164: out<=1;
   58165: out<=1;
   58166: out<=0;
   58167: out<=0;
   58168: out<=0;
   58169: out<=0;
   58170: out<=0;
   58171: out<=0;
   58172: out<=1;
   58173: out<=0;
   58174: out<=0;
   58175: out<=1;
   58176: out<=1;
   58177: out<=0;
   58178: out<=0;
   58179: out<=1;
   58180: out<=0;
   58181: out<=0;
   58182: out<=0;
   58183: out<=0;
   58184: out<=0;
   58185: out<=0;
   58186: out<=1;
   58187: out<=1;
   58188: out<=1;
   58189: out<=0;
   58190: out<=1;
   58191: out<=0;
   58192: out<=1;
   58193: out<=1;
   58194: out<=1;
   58195: out<=1;
   58196: out<=1;
   58197: out<=0;
   58198: out<=0;
   58199: out<=1;
   58200: out<=1;
   58201: out<=0;
   58202: out<=1;
   58203: out<=0;
   58204: out<=1;
   58205: out<=1;
   58206: out<=0;
   58207: out<=0;
   58208: out<=1;
   58209: out<=1;
   58210: out<=0;
   58211: out<=0;
   58212: out<=1;
   58213: out<=0;
   58214: out<=1;
   58215: out<=0;
   58216: out<=0;
   58217: out<=1;
   58218: out<=1;
   58219: out<=0;
   58220: out<=0;
   58221: out<=0;
   58222: out<=0;
   58223: out<=0;
   58224: out<=1;
   58225: out<=0;
   58226: out<=1;
   58227: out<=0;
   58228: out<=0;
   58229: out<=0;
   58230: out<=1;
   58231: out<=1;
   58232: out<=1;
   58233: out<=1;
   58234: out<=1;
   58235: out<=1;
   58236: out<=0;
   58237: out<=1;
   58238: out<=1;
   58239: out<=0;
   58240: out<=0;
   58241: out<=1;
   58242: out<=1;
   58243: out<=0;
   58244: out<=1;
   58245: out<=1;
   58246: out<=1;
   58247: out<=1;
   58248: out<=1;
   58249: out<=1;
   58250: out<=0;
   58251: out<=0;
   58252: out<=0;
   58253: out<=1;
   58254: out<=0;
   58255: out<=1;
   58256: out<=0;
   58257: out<=0;
   58258: out<=0;
   58259: out<=0;
   58260: out<=0;
   58261: out<=1;
   58262: out<=1;
   58263: out<=0;
   58264: out<=0;
   58265: out<=1;
   58266: out<=0;
   58267: out<=1;
   58268: out<=0;
   58269: out<=0;
   58270: out<=1;
   58271: out<=1;
   58272: out<=1;
   58273: out<=1;
   58274: out<=0;
   58275: out<=0;
   58276: out<=1;
   58277: out<=0;
   58278: out<=1;
   58279: out<=0;
   58280: out<=0;
   58281: out<=1;
   58282: out<=1;
   58283: out<=0;
   58284: out<=0;
   58285: out<=0;
   58286: out<=0;
   58287: out<=0;
   58288: out<=1;
   58289: out<=0;
   58290: out<=1;
   58291: out<=0;
   58292: out<=0;
   58293: out<=0;
   58294: out<=1;
   58295: out<=1;
   58296: out<=1;
   58297: out<=1;
   58298: out<=1;
   58299: out<=1;
   58300: out<=0;
   58301: out<=1;
   58302: out<=1;
   58303: out<=0;
   58304: out<=1;
   58305: out<=0;
   58306: out<=0;
   58307: out<=1;
   58308: out<=0;
   58309: out<=0;
   58310: out<=0;
   58311: out<=0;
   58312: out<=0;
   58313: out<=0;
   58314: out<=1;
   58315: out<=1;
   58316: out<=1;
   58317: out<=0;
   58318: out<=1;
   58319: out<=0;
   58320: out<=0;
   58321: out<=0;
   58322: out<=0;
   58323: out<=0;
   58324: out<=0;
   58325: out<=1;
   58326: out<=1;
   58327: out<=0;
   58328: out<=0;
   58329: out<=1;
   58330: out<=0;
   58331: out<=1;
   58332: out<=0;
   58333: out<=0;
   58334: out<=1;
   58335: out<=1;
   58336: out<=1;
   58337: out<=1;
   58338: out<=0;
   58339: out<=0;
   58340: out<=1;
   58341: out<=0;
   58342: out<=1;
   58343: out<=0;
   58344: out<=0;
   58345: out<=1;
   58346: out<=1;
   58347: out<=0;
   58348: out<=0;
   58349: out<=0;
   58350: out<=0;
   58351: out<=0;
   58352: out<=0;
   58353: out<=1;
   58354: out<=0;
   58355: out<=1;
   58356: out<=1;
   58357: out<=1;
   58358: out<=0;
   58359: out<=0;
   58360: out<=0;
   58361: out<=0;
   58362: out<=0;
   58363: out<=0;
   58364: out<=1;
   58365: out<=0;
   58366: out<=0;
   58367: out<=1;
   58368: out<=1;
   58369: out<=1;
   58370: out<=0;
   58371: out<=0;
   58372: out<=0;
   58373: out<=1;
   58374: out<=0;
   58375: out<=1;
   58376: out<=1;
   58377: out<=0;
   58378: out<=0;
   58379: out<=1;
   58380: out<=0;
   58381: out<=0;
   58382: out<=0;
   58383: out<=0;
   58384: out<=0;
   58385: out<=1;
   58386: out<=0;
   58387: out<=1;
   58388: out<=0;
   58389: out<=0;
   58390: out<=1;
   58391: out<=1;
   58392: out<=1;
   58393: out<=1;
   58394: out<=1;
   58395: out<=1;
   58396: out<=1;
   58397: out<=0;
   58398: out<=0;
   58399: out<=1;
   58400: out<=1;
   58401: out<=0;
   58402: out<=0;
   58403: out<=1;
   58404: out<=1;
   58405: out<=1;
   58406: out<=1;
   58407: out<=1;
   58408: out<=1;
   58409: out<=1;
   58410: out<=0;
   58411: out<=0;
   58412: out<=1;
   58413: out<=0;
   58414: out<=1;
   58415: out<=0;
   58416: out<=0;
   58417: out<=0;
   58418: out<=0;
   58419: out<=0;
   58420: out<=1;
   58421: out<=0;
   58422: out<=0;
   58423: out<=1;
   58424: out<=1;
   58425: out<=0;
   58426: out<=1;
   58427: out<=0;
   58428: out<=0;
   58429: out<=0;
   58430: out<=1;
   58431: out<=1;
   58432: out<=1;
   58433: out<=1;
   58434: out<=0;
   58435: out<=0;
   58436: out<=0;
   58437: out<=1;
   58438: out<=0;
   58439: out<=1;
   58440: out<=1;
   58441: out<=0;
   58442: out<=0;
   58443: out<=1;
   58444: out<=0;
   58445: out<=0;
   58446: out<=0;
   58447: out<=0;
   58448: out<=1;
   58449: out<=0;
   58450: out<=1;
   58451: out<=0;
   58452: out<=1;
   58453: out<=1;
   58454: out<=0;
   58455: out<=0;
   58456: out<=0;
   58457: out<=0;
   58458: out<=0;
   58459: out<=0;
   58460: out<=0;
   58461: out<=1;
   58462: out<=1;
   58463: out<=0;
   58464: out<=0;
   58465: out<=1;
   58466: out<=1;
   58467: out<=0;
   58468: out<=0;
   58469: out<=0;
   58470: out<=0;
   58471: out<=0;
   58472: out<=0;
   58473: out<=0;
   58474: out<=1;
   58475: out<=1;
   58476: out<=0;
   58477: out<=1;
   58478: out<=0;
   58479: out<=1;
   58480: out<=0;
   58481: out<=0;
   58482: out<=0;
   58483: out<=0;
   58484: out<=1;
   58485: out<=0;
   58486: out<=0;
   58487: out<=1;
   58488: out<=1;
   58489: out<=0;
   58490: out<=1;
   58491: out<=0;
   58492: out<=0;
   58493: out<=0;
   58494: out<=1;
   58495: out<=1;
   58496: out<=1;
   58497: out<=1;
   58498: out<=0;
   58499: out<=0;
   58500: out<=0;
   58501: out<=1;
   58502: out<=0;
   58503: out<=1;
   58504: out<=1;
   58505: out<=0;
   58506: out<=0;
   58507: out<=1;
   58508: out<=0;
   58509: out<=0;
   58510: out<=0;
   58511: out<=0;
   58512: out<=1;
   58513: out<=0;
   58514: out<=1;
   58515: out<=0;
   58516: out<=1;
   58517: out<=1;
   58518: out<=0;
   58519: out<=0;
   58520: out<=0;
   58521: out<=0;
   58522: out<=0;
   58523: out<=0;
   58524: out<=0;
   58525: out<=1;
   58526: out<=1;
   58527: out<=0;
   58528: out<=1;
   58529: out<=0;
   58530: out<=0;
   58531: out<=1;
   58532: out<=1;
   58533: out<=1;
   58534: out<=1;
   58535: out<=1;
   58536: out<=1;
   58537: out<=1;
   58538: out<=0;
   58539: out<=0;
   58540: out<=1;
   58541: out<=0;
   58542: out<=1;
   58543: out<=0;
   58544: out<=1;
   58545: out<=1;
   58546: out<=1;
   58547: out<=1;
   58548: out<=0;
   58549: out<=1;
   58550: out<=1;
   58551: out<=0;
   58552: out<=0;
   58553: out<=1;
   58554: out<=0;
   58555: out<=1;
   58556: out<=1;
   58557: out<=1;
   58558: out<=0;
   58559: out<=0;
   58560: out<=1;
   58561: out<=1;
   58562: out<=0;
   58563: out<=0;
   58564: out<=0;
   58565: out<=1;
   58566: out<=0;
   58567: out<=1;
   58568: out<=1;
   58569: out<=0;
   58570: out<=0;
   58571: out<=1;
   58572: out<=0;
   58573: out<=0;
   58574: out<=0;
   58575: out<=0;
   58576: out<=0;
   58577: out<=1;
   58578: out<=0;
   58579: out<=1;
   58580: out<=0;
   58581: out<=0;
   58582: out<=1;
   58583: out<=1;
   58584: out<=1;
   58585: out<=1;
   58586: out<=1;
   58587: out<=1;
   58588: out<=1;
   58589: out<=0;
   58590: out<=0;
   58591: out<=1;
   58592: out<=0;
   58593: out<=1;
   58594: out<=1;
   58595: out<=0;
   58596: out<=0;
   58597: out<=0;
   58598: out<=0;
   58599: out<=0;
   58600: out<=0;
   58601: out<=0;
   58602: out<=1;
   58603: out<=1;
   58604: out<=0;
   58605: out<=1;
   58606: out<=0;
   58607: out<=1;
   58608: out<=1;
   58609: out<=1;
   58610: out<=1;
   58611: out<=1;
   58612: out<=0;
   58613: out<=1;
   58614: out<=1;
   58615: out<=0;
   58616: out<=0;
   58617: out<=1;
   58618: out<=0;
   58619: out<=1;
   58620: out<=1;
   58621: out<=1;
   58622: out<=0;
   58623: out<=0;
   58624: out<=1;
   58625: out<=0;
   58626: out<=1;
   58627: out<=0;
   58628: out<=1;
   58629: out<=1;
   58630: out<=0;
   58631: out<=0;
   58632: out<=0;
   58633: out<=0;
   58634: out<=0;
   58635: out<=0;
   58636: out<=0;
   58637: out<=1;
   58638: out<=1;
   58639: out<=0;
   58640: out<=1;
   58641: out<=1;
   58642: out<=0;
   58643: out<=0;
   58644: out<=0;
   58645: out<=1;
   58646: out<=0;
   58647: out<=1;
   58648: out<=1;
   58649: out<=0;
   58650: out<=0;
   58651: out<=1;
   58652: out<=0;
   58653: out<=0;
   58654: out<=0;
   58655: out<=0;
   58656: out<=0;
   58657: out<=0;
   58658: out<=0;
   58659: out<=0;
   58660: out<=1;
   58661: out<=0;
   58662: out<=0;
   58663: out<=1;
   58664: out<=1;
   58665: out<=0;
   58666: out<=1;
   58667: out<=0;
   58668: out<=0;
   58669: out<=0;
   58670: out<=1;
   58671: out<=1;
   58672: out<=0;
   58673: out<=1;
   58674: out<=1;
   58675: out<=0;
   58676: out<=0;
   58677: out<=0;
   58678: out<=0;
   58679: out<=0;
   58680: out<=0;
   58681: out<=0;
   58682: out<=1;
   58683: out<=1;
   58684: out<=0;
   58685: out<=1;
   58686: out<=0;
   58687: out<=1;
   58688: out<=0;
   58689: out<=1;
   58690: out<=0;
   58691: out<=1;
   58692: out<=0;
   58693: out<=0;
   58694: out<=1;
   58695: out<=1;
   58696: out<=1;
   58697: out<=1;
   58698: out<=1;
   58699: out<=1;
   58700: out<=1;
   58701: out<=0;
   58702: out<=0;
   58703: out<=1;
   58704: out<=1;
   58705: out<=1;
   58706: out<=0;
   58707: out<=0;
   58708: out<=0;
   58709: out<=1;
   58710: out<=0;
   58711: out<=1;
   58712: out<=1;
   58713: out<=0;
   58714: out<=0;
   58715: out<=1;
   58716: out<=0;
   58717: out<=0;
   58718: out<=0;
   58719: out<=0;
   58720: out<=0;
   58721: out<=0;
   58722: out<=0;
   58723: out<=0;
   58724: out<=1;
   58725: out<=0;
   58726: out<=0;
   58727: out<=1;
   58728: out<=1;
   58729: out<=0;
   58730: out<=1;
   58731: out<=0;
   58732: out<=0;
   58733: out<=0;
   58734: out<=1;
   58735: out<=1;
   58736: out<=1;
   58737: out<=0;
   58738: out<=0;
   58739: out<=1;
   58740: out<=1;
   58741: out<=1;
   58742: out<=1;
   58743: out<=1;
   58744: out<=1;
   58745: out<=1;
   58746: out<=0;
   58747: out<=0;
   58748: out<=1;
   58749: out<=0;
   58750: out<=1;
   58751: out<=0;
   58752: out<=0;
   58753: out<=1;
   58754: out<=0;
   58755: out<=1;
   58756: out<=0;
   58757: out<=0;
   58758: out<=1;
   58759: out<=1;
   58760: out<=1;
   58761: out<=1;
   58762: out<=1;
   58763: out<=1;
   58764: out<=1;
   58765: out<=0;
   58766: out<=0;
   58767: out<=1;
   58768: out<=1;
   58769: out<=1;
   58770: out<=0;
   58771: out<=0;
   58772: out<=0;
   58773: out<=1;
   58774: out<=0;
   58775: out<=1;
   58776: out<=1;
   58777: out<=0;
   58778: out<=0;
   58779: out<=1;
   58780: out<=0;
   58781: out<=0;
   58782: out<=0;
   58783: out<=0;
   58784: out<=1;
   58785: out<=1;
   58786: out<=1;
   58787: out<=1;
   58788: out<=0;
   58789: out<=1;
   58790: out<=1;
   58791: out<=0;
   58792: out<=0;
   58793: out<=1;
   58794: out<=0;
   58795: out<=1;
   58796: out<=1;
   58797: out<=1;
   58798: out<=0;
   58799: out<=0;
   58800: out<=0;
   58801: out<=1;
   58802: out<=1;
   58803: out<=0;
   58804: out<=0;
   58805: out<=0;
   58806: out<=0;
   58807: out<=0;
   58808: out<=0;
   58809: out<=0;
   58810: out<=1;
   58811: out<=1;
   58812: out<=0;
   58813: out<=1;
   58814: out<=0;
   58815: out<=1;
   58816: out<=1;
   58817: out<=0;
   58818: out<=1;
   58819: out<=0;
   58820: out<=1;
   58821: out<=1;
   58822: out<=0;
   58823: out<=0;
   58824: out<=0;
   58825: out<=0;
   58826: out<=0;
   58827: out<=0;
   58828: out<=0;
   58829: out<=1;
   58830: out<=1;
   58831: out<=0;
   58832: out<=1;
   58833: out<=1;
   58834: out<=0;
   58835: out<=0;
   58836: out<=0;
   58837: out<=1;
   58838: out<=0;
   58839: out<=1;
   58840: out<=1;
   58841: out<=0;
   58842: out<=0;
   58843: out<=1;
   58844: out<=0;
   58845: out<=0;
   58846: out<=0;
   58847: out<=0;
   58848: out<=1;
   58849: out<=1;
   58850: out<=1;
   58851: out<=1;
   58852: out<=0;
   58853: out<=1;
   58854: out<=1;
   58855: out<=0;
   58856: out<=0;
   58857: out<=1;
   58858: out<=0;
   58859: out<=1;
   58860: out<=1;
   58861: out<=1;
   58862: out<=0;
   58863: out<=0;
   58864: out<=1;
   58865: out<=0;
   58866: out<=0;
   58867: out<=1;
   58868: out<=1;
   58869: out<=1;
   58870: out<=1;
   58871: out<=1;
   58872: out<=1;
   58873: out<=1;
   58874: out<=0;
   58875: out<=0;
   58876: out<=1;
   58877: out<=0;
   58878: out<=1;
   58879: out<=0;
   58880: out<=1;
   58881: out<=0;
   58882: out<=0;
   58883: out<=1;
   58884: out<=1;
   58885: out<=1;
   58886: out<=1;
   58887: out<=1;
   58888: out<=1;
   58889: out<=1;
   58890: out<=0;
   58891: out<=0;
   58892: out<=1;
   58893: out<=0;
   58894: out<=1;
   58895: out<=0;
   58896: out<=1;
   58897: out<=1;
   58898: out<=1;
   58899: out<=1;
   58900: out<=0;
   58901: out<=1;
   58902: out<=1;
   58903: out<=0;
   58904: out<=0;
   58905: out<=1;
   58906: out<=0;
   58907: out<=1;
   58908: out<=1;
   58909: out<=1;
   58910: out<=0;
   58911: out<=0;
   58912: out<=1;
   58913: out<=1;
   58914: out<=0;
   58915: out<=0;
   58916: out<=0;
   58917: out<=1;
   58918: out<=0;
   58919: out<=1;
   58920: out<=1;
   58921: out<=0;
   58922: out<=0;
   58923: out<=1;
   58924: out<=0;
   58925: out<=0;
   58926: out<=0;
   58927: out<=0;
   58928: out<=1;
   58929: out<=0;
   58930: out<=1;
   58931: out<=0;
   58932: out<=1;
   58933: out<=1;
   58934: out<=0;
   58935: out<=0;
   58936: out<=0;
   58937: out<=0;
   58938: out<=0;
   58939: out<=0;
   58940: out<=0;
   58941: out<=1;
   58942: out<=1;
   58943: out<=0;
   58944: out<=0;
   58945: out<=1;
   58946: out<=1;
   58947: out<=0;
   58948: out<=0;
   58949: out<=0;
   58950: out<=0;
   58951: out<=0;
   58952: out<=0;
   58953: out<=0;
   58954: out<=1;
   58955: out<=1;
   58956: out<=0;
   58957: out<=1;
   58958: out<=0;
   58959: out<=1;
   58960: out<=1;
   58961: out<=1;
   58962: out<=1;
   58963: out<=1;
   58964: out<=0;
   58965: out<=1;
   58966: out<=1;
   58967: out<=0;
   58968: out<=0;
   58969: out<=1;
   58970: out<=0;
   58971: out<=1;
   58972: out<=1;
   58973: out<=1;
   58974: out<=0;
   58975: out<=0;
   58976: out<=1;
   58977: out<=1;
   58978: out<=0;
   58979: out<=0;
   58980: out<=0;
   58981: out<=1;
   58982: out<=0;
   58983: out<=1;
   58984: out<=1;
   58985: out<=0;
   58986: out<=0;
   58987: out<=1;
   58988: out<=0;
   58989: out<=0;
   58990: out<=0;
   58991: out<=0;
   58992: out<=0;
   58993: out<=1;
   58994: out<=0;
   58995: out<=1;
   58996: out<=0;
   58997: out<=0;
   58998: out<=1;
   58999: out<=1;
   59000: out<=1;
   59001: out<=1;
   59002: out<=1;
   59003: out<=1;
   59004: out<=1;
   59005: out<=0;
   59006: out<=0;
   59007: out<=1;
   59008: out<=1;
   59009: out<=0;
   59010: out<=0;
   59011: out<=1;
   59012: out<=1;
   59013: out<=1;
   59014: out<=1;
   59015: out<=1;
   59016: out<=1;
   59017: out<=1;
   59018: out<=0;
   59019: out<=0;
   59020: out<=1;
   59021: out<=0;
   59022: out<=1;
   59023: out<=0;
   59024: out<=0;
   59025: out<=0;
   59026: out<=0;
   59027: out<=0;
   59028: out<=1;
   59029: out<=0;
   59030: out<=0;
   59031: out<=1;
   59032: out<=1;
   59033: out<=0;
   59034: out<=1;
   59035: out<=0;
   59036: out<=0;
   59037: out<=0;
   59038: out<=1;
   59039: out<=1;
   59040: out<=1;
   59041: out<=1;
   59042: out<=0;
   59043: out<=0;
   59044: out<=0;
   59045: out<=1;
   59046: out<=0;
   59047: out<=1;
   59048: out<=1;
   59049: out<=0;
   59050: out<=0;
   59051: out<=1;
   59052: out<=0;
   59053: out<=0;
   59054: out<=0;
   59055: out<=0;
   59056: out<=0;
   59057: out<=1;
   59058: out<=0;
   59059: out<=1;
   59060: out<=0;
   59061: out<=0;
   59062: out<=1;
   59063: out<=1;
   59064: out<=1;
   59065: out<=1;
   59066: out<=1;
   59067: out<=1;
   59068: out<=1;
   59069: out<=0;
   59070: out<=0;
   59071: out<=1;
   59072: out<=0;
   59073: out<=1;
   59074: out<=1;
   59075: out<=0;
   59076: out<=0;
   59077: out<=0;
   59078: out<=0;
   59079: out<=0;
   59080: out<=0;
   59081: out<=0;
   59082: out<=1;
   59083: out<=1;
   59084: out<=0;
   59085: out<=1;
   59086: out<=0;
   59087: out<=1;
   59088: out<=0;
   59089: out<=0;
   59090: out<=0;
   59091: out<=0;
   59092: out<=1;
   59093: out<=0;
   59094: out<=0;
   59095: out<=1;
   59096: out<=1;
   59097: out<=0;
   59098: out<=1;
   59099: out<=0;
   59100: out<=0;
   59101: out<=0;
   59102: out<=1;
   59103: out<=1;
   59104: out<=1;
   59105: out<=1;
   59106: out<=0;
   59107: out<=0;
   59108: out<=0;
   59109: out<=1;
   59110: out<=0;
   59111: out<=1;
   59112: out<=1;
   59113: out<=0;
   59114: out<=0;
   59115: out<=1;
   59116: out<=0;
   59117: out<=0;
   59118: out<=0;
   59119: out<=0;
   59120: out<=1;
   59121: out<=0;
   59122: out<=1;
   59123: out<=0;
   59124: out<=1;
   59125: out<=1;
   59126: out<=0;
   59127: out<=0;
   59128: out<=0;
   59129: out<=0;
   59130: out<=0;
   59131: out<=0;
   59132: out<=0;
   59133: out<=1;
   59134: out<=1;
   59135: out<=0;
   59136: out<=1;
   59137: out<=1;
   59138: out<=1;
   59139: out<=1;
   59140: out<=0;
   59141: out<=1;
   59142: out<=1;
   59143: out<=0;
   59144: out<=0;
   59145: out<=1;
   59146: out<=0;
   59147: out<=1;
   59148: out<=1;
   59149: out<=1;
   59150: out<=0;
   59151: out<=0;
   59152: out<=0;
   59153: out<=1;
   59154: out<=1;
   59155: out<=0;
   59156: out<=0;
   59157: out<=0;
   59158: out<=0;
   59159: out<=0;
   59160: out<=0;
   59161: out<=0;
   59162: out<=1;
   59163: out<=1;
   59164: out<=0;
   59165: out<=1;
   59166: out<=0;
   59167: out<=1;
   59168: out<=0;
   59169: out<=1;
   59170: out<=0;
   59171: out<=1;
   59172: out<=0;
   59173: out<=0;
   59174: out<=1;
   59175: out<=1;
   59176: out<=1;
   59177: out<=1;
   59178: out<=1;
   59179: out<=1;
   59180: out<=1;
   59181: out<=0;
   59182: out<=0;
   59183: out<=1;
   59184: out<=1;
   59185: out<=1;
   59186: out<=0;
   59187: out<=0;
   59188: out<=0;
   59189: out<=1;
   59190: out<=0;
   59191: out<=1;
   59192: out<=1;
   59193: out<=0;
   59194: out<=0;
   59195: out<=1;
   59196: out<=0;
   59197: out<=0;
   59198: out<=0;
   59199: out<=0;
   59200: out<=1;
   59201: out<=1;
   59202: out<=1;
   59203: out<=1;
   59204: out<=0;
   59205: out<=1;
   59206: out<=1;
   59207: out<=0;
   59208: out<=0;
   59209: out<=1;
   59210: out<=0;
   59211: out<=1;
   59212: out<=1;
   59213: out<=1;
   59214: out<=0;
   59215: out<=0;
   59216: out<=1;
   59217: out<=0;
   59218: out<=0;
   59219: out<=1;
   59220: out<=1;
   59221: out<=1;
   59222: out<=1;
   59223: out<=1;
   59224: out<=1;
   59225: out<=1;
   59226: out<=0;
   59227: out<=0;
   59228: out<=1;
   59229: out<=0;
   59230: out<=1;
   59231: out<=0;
   59232: out<=1;
   59233: out<=0;
   59234: out<=1;
   59235: out<=0;
   59236: out<=1;
   59237: out<=1;
   59238: out<=0;
   59239: out<=0;
   59240: out<=0;
   59241: out<=0;
   59242: out<=0;
   59243: out<=0;
   59244: out<=0;
   59245: out<=1;
   59246: out<=1;
   59247: out<=0;
   59248: out<=1;
   59249: out<=1;
   59250: out<=0;
   59251: out<=0;
   59252: out<=0;
   59253: out<=1;
   59254: out<=0;
   59255: out<=1;
   59256: out<=1;
   59257: out<=0;
   59258: out<=0;
   59259: out<=1;
   59260: out<=0;
   59261: out<=0;
   59262: out<=0;
   59263: out<=0;
   59264: out<=0;
   59265: out<=0;
   59266: out<=0;
   59267: out<=0;
   59268: out<=1;
   59269: out<=0;
   59270: out<=0;
   59271: out<=1;
   59272: out<=1;
   59273: out<=0;
   59274: out<=1;
   59275: out<=0;
   59276: out<=0;
   59277: out<=0;
   59278: out<=1;
   59279: out<=1;
   59280: out<=0;
   59281: out<=1;
   59282: out<=1;
   59283: out<=0;
   59284: out<=0;
   59285: out<=0;
   59286: out<=0;
   59287: out<=0;
   59288: out<=0;
   59289: out<=0;
   59290: out<=1;
   59291: out<=1;
   59292: out<=0;
   59293: out<=1;
   59294: out<=0;
   59295: out<=1;
   59296: out<=1;
   59297: out<=0;
   59298: out<=1;
   59299: out<=0;
   59300: out<=1;
   59301: out<=1;
   59302: out<=0;
   59303: out<=0;
   59304: out<=0;
   59305: out<=0;
   59306: out<=0;
   59307: out<=0;
   59308: out<=0;
   59309: out<=1;
   59310: out<=1;
   59311: out<=0;
   59312: out<=1;
   59313: out<=1;
   59314: out<=0;
   59315: out<=0;
   59316: out<=0;
   59317: out<=1;
   59318: out<=0;
   59319: out<=1;
   59320: out<=1;
   59321: out<=0;
   59322: out<=0;
   59323: out<=1;
   59324: out<=0;
   59325: out<=0;
   59326: out<=0;
   59327: out<=0;
   59328: out<=0;
   59329: out<=0;
   59330: out<=0;
   59331: out<=0;
   59332: out<=1;
   59333: out<=0;
   59334: out<=0;
   59335: out<=1;
   59336: out<=1;
   59337: out<=0;
   59338: out<=1;
   59339: out<=0;
   59340: out<=0;
   59341: out<=0;
   59342: out<=1;
   59343: out<=1;
   59344: out<=1;
   59345: out<=0;
   59346: out<=0;
   59347: out<=1;
   59348: out<=1;
   59349: out<=1;
   59350: out<=1;
   59351: out<=1;
   59352: out<=1;
   59353: out<=1;
   59354: out<=0;
   59355: out<=0;
   59356: out<=1;
   59357: out<=0;
   59358: out<=1;
   59359: out<=0;
   59360: out<=0;
   59361: out<=1;
   59362: out<=0;
   59363: out<=1;
   59364: out<=0;
   59365: out<=0;
   59366: out<=1;
   59367: out<=1;
   59368: out<=1;
   59369: out<=1;
   59370: out<=1;
   59371: out<=1;
   59372: out<=1;
   59373: out<=0;
   59374: out<=0;
   59375: out<=1;
   59376: out<=1;
   59377: out<=1;
   59378: out<=0;
   59379: out<=0;
   59380: out<=0;
   59381: out<=1;
   59382: out<=0;
   59383: out<=1;
   59384: out<=1;
   59385: out<=0;
   59386: out<=0;
   59387: out<=1;
   59388: out<=0;
   59389: out<=0;
   59390: out<=0;
   59391: out<=0;
   59392: out<=1;
   59393: out<=1;
   59394: out<=1;
   59395: out<=1;
   59396: out<=0;
   59397: out<=1;
   59398: out<=1;
   59399: out<=0;
   59400: out<=1;
   59401: out<=0;
   59402: out<=1;
   59403: out<=0;
   59404: out<=0;
   59405: out<=0;
   59406: out<=1;
   59407: out<=1;
   59408: out<=0;
   59409: out<=1;
   59410: out<=1;
   59411: out<=0;
   59412: out<=0;
   59413: out<=0;
   59414: out<=0;
   59415: out<=0;
   59416: out<=1;
   59417: out<=1;
   59418: out<=0;
   59419: out<=0;
   59420: out<=1;
   59421: out<=0;
   59422: out<=1;
   59423: out<=0;
   59424: out<=1;
   59425: out<=0;
   59426: out<=1;
   59427: out<=0;
   59428: out<=1;
   59429: out<=1;
   59430: out<=0;
   59431: out<=0;
   59432: out<=1;
   59433: out<=1;
   59434: out<=1;
   59435: out<=1;
   59436: out<=1;
   59437: out<=0;
   59438: out<=0;
   59439: out<=1;
   59440: out<=0;
   59441: out<=0;
   59442: out<=1;
   59443: out<=1;
   59444: out<=1;
   59445: out<=0;
   59446: out<=1;
   59447: out<=0;
   59448: out<=1;
   59449: out<=0;
   59450: out<=0;
   59451: out<=1;
   59452: out<=0;
   59453: out<=0;
   59454: out<=0;
   59455: out<=0;
   59456: out<=1;
   59457: out<=1;
   59458: out<=1;
   59459: out<=1;
   59460: out<=0;
   59461: out<=1;
   59462: out<=1;
   59463: out<=0;
   59464: out<=1;
   59465: out<=0;
   59466: out<=1;
   59467: out<=0;
   59468: out<=0;
   59469: out<=0;
   59470: out<=1;
   59471: out<=1;
   59472: out<=1;
   59473: out<=0;
   59474: out<=0;
   59475: out<=1;
   59476: out<=1;
   59477: out<=1;
   59478: out<=1;
   59479: out<=1;
   59480: out<=0;
   59481: out<=0;
   59482: out<=1;
   59483: out<=1;
   59484: out<=0;
   59485: out<=1;
   59486: out<=0;
   59487: out<=1;
   59488: out<=0;
   59489: out<=1;
   59490: out<=0;
   59491: out<=1;
   59492: out<=0;
   59493: out<=0;
   59494: out<=1;
   59495: out<=1;
   59496: out<=0;
   59497: out<=0;
   59498: out<=0;
   59499: out<=0;
   59500: out<=0;
   59501: out<=1;
   59502: out<=1;
   59503: out<=0;
   59504: out<=0;
   59505: out<=0;
   59506: out<=1;
   59507: out<=1;
   59508: out<=1;
   59509: out<=0;
   59510: out<=1;
   59511: out<=0;
   59512: out<=1;
   59513: out<=0;
   59514: out<=0;
   59515: out<=1;
   59516: out<=0;
   59517: out<=0;
   59518: out<=0;
   59519: out<=0;
   59520: out<=0;
   59521: out<=0;
   59522: out<=0;
   59523: out<=0;
   59524: out<=1;
   59525: out<=0;
   59526: out<=0;
   59527: out<=1;
   59528: out<=0;
   59529: out<=1;
   59530: out<=0;
   59531: out<=1;
   59532: out<=1;
   59533: out<=1;
   59534: out<=0;
   59535: out<=0;
   59536: out<=0;
   59537: out<=1;
   59538: out<=1;
   59539: out<=0;
   59540: out<=0;
   59541: out<=0;
   59542: out<=0;
   59543: out<=0;
   59544: out<=1;
   59545: out<=1;
   59546: out<=0;
   59547: out<=0;
   59548: out<=1;
   59549: out<=0;
   59550: out<=1;
   59551: out<=0;
   59552: out<=0;
   59553: out<=1;
   59554: out<=0;
   59555: out<=1;
   59556: out<=0;
   59557: out<=0;
   59558: out<=1;
   59559: out<=1;
   59560: out<=0;
   59561: out<=0;
   59562: out<=0;
   59563: out<=0;
   59564: out<=0;
   59565: out<=1;
   59566: out<=1;
   59567: out<=0;
   59568: out<=0;
   59569: out<=0;
   59570: out<=1;
   59571: out<=1;
   59572: out<=1;
   59573: out<=0;
   59574: out<=1;
   59575: out<=0;
   59576: out<=1;
   59577: out<=0;
   59578: out<=0;
   59579: out<=1;
   59580: out<=0;
   59581: out<=0;
   59582: out<=0;
   59583: out<=0;
   59584: out<=0;
   59585: out<=0;
   59586: out<=0;
   59587: out<=0;
   59588: out<=1;
   59589: out<=0;
   59590: out<=0;
   59591: out<=1;
   59592: out<=0;
   59593: out<=1;
   59594: out<=0;
   59595: out<=1;
   59596: out<=1;
   59597: out<=1;
   59598: out<=0;
   59599: out<=0;
   59600: out<=1;
   59601: out<=0;
   59602: out<=0;
   59603: out<=1;
   59604: out<=1;
   59605: out<=1;
   59606: out<=1;
   59607: out<=1;
   59608: out<=0;
   59609: out<=0;
   59610: out<=1;
   59611: out<=1;
   59612: out<=0;
   59613: out<=1;
   59614: out<=0;
   59615: out<=1;
   59616: out<=1;
   59617: out<=0;
   59618: out<=1;
   59619: out<=0;
   59620: out<=1;
   59621: out<=1;
   59622: out<=0;
   59623: out<=0;
   59624: out<=1;
   59625: out<=1;
   59626: out<=1;
   59627: out<=1;
   59628: out<=1;
   59629: out<=0;
   59630: out<=0;
   59631: out<=1;
   59632: out<=0;
   59633: out<=0;
   59634: out<=1;
   59635: out<=1;
   59636: out<=1;
   59637: out<=0;
   59638: out<=1;
   59639: out<=0;
   59640: out<=1;
   59641: out<=0;
   59642: out<=0;
   59643: out<=1;
   59644: out<=0;
   59645: out<=0;
   59646: out<=0;
   59647: out<=0;
   59648: out<=1;
   59649: out<=0;
   59650: out<=0;
   59651: out<=1;
   59652: out<=1;
   59653: out<=1;
   59654: out<=1;
   59655: out<=1;
   59656: out<=0;
   59657: out<=0;
   59658: out<=1;
   59659: out<=1;
   59660: out<=0;
   59661: out<=1;
   59662: out<=0;
   59663: out<=1;
   59664: out<=1;
   59665: out<=1;
   59666: out<=1;
   59667: out<=1;
   59668: out<=0;
   59669: out<=1;
   59670: out<=1;
   59671: out<=0;
   59672: out<=1;
   59673: out<=0;
   59674: out<=1;
   59675: out<=0;
   59676: out<=0;
   59677: out<=0;
   59678: out<=1;
   59679: out<=1;
   59680: out<=0;
   59681: out<=0;
   59682: out<=1;
   59683: out<=1;
   59684: out<=1;
   59685: out<=0;
   59686: out<=1;
   59687: out<=0;
   59688: out<=1;
   59689: out<=0;
   59690: out<=0;
   59691: out<=1;
   59692: out<=0;
   59693: out<=0;
   59694: out<=0;
   59695: out<=0;
   59696: out<=0;
   59697: out<=1;
   59698: out<=0;
   59699: out<=1;
   59700: out<=0;
   59701: out<=0;
   59702: out<=1;
   59703: out<=1;
   59704: out<=0;
   59705: out<=0;
   59706: out<=0;
   59707: out<=0;
   59708: out<=0;
   59709: out<=1;
   59710: out<=1;
   59711: out<=0;
   59712: out<=0;
   59713: out<=1;
   59714: out<=1;
   59715: out<=0;
   59716: out<=0;
   59717: out<=0;
   59718: out<=0;
   59719: out<=0;
   59720: out<=1;
   59721: out<=1;
   59722: out<=0;
   59723: out<=0;
   59724: out<=1;
   59725: out<=0;
   59726: out<=1;
   59727: out<=0;
   59728: out<=1;
   59729: out<=1;
   59730: out<=1;
   59731: out<=1;
   59732: out<=0;
   59733: out<=1;
   59734: out<=1;
   59735: out<=0;
   59736: out<=1;
   59737: out<=0;
   59738: out<=1;
   59739: out<=0;
   59740: out<=0;
   59741: out<=0;
   59742: out<=1;
   59743: out<=1;
   59744: out<=0;
   59745: out<=0;
   59746: out<=1;
   59747: out<=1;
   59748: out<=1;
   59749: out<=0;
   59750: out<=1;
   59751: out<=0;
   59752: out<=1;
   59753: out<=0;
   59754: out<=0;
   59755: out<=1;
   59756: out<=0;
   59757: out<=0;
   59758: out<=0;
   59759: out<=0;
   59760: out<=1;
   59761: out<=0;
   59762: out<=1;
   59763: out<=0;
   59764: out<=1;
   59765: out<=1;
   59766: out<=0;
   59767: out<=0;
   59768: out<=1;
   59769: out<=1;
   59770: out<=1;
   59771: out<=1;
   59772: out<=1;
   59773: out<=0;
   59774: out<=0;
   59775: out<=1;
   59776: out<=1;
   59777: out<=0;
   59778: out<=0;
   59779: out<=1;
   59780: out<=1;
   59781: out<=1;
   59782: out<=1;
   59783: out<=1;
   59784: out<=0;
   59785: out<=0;
   59786: out<=1;
   59787: out<=1;
   59788: out<=0;
   59789: out<=1;
   59790: out<=0;
   59791: out<=1;
   59792: out<=0;
   59793: out<=0;
   59794: out<=0;
   59795: out<=0;
   59796: out<=1;
   59797: out<=0;
   59798: out<=0;
   59799: out<=1;
   59800: out<=0;
   59801: out<=1;
   59802: out<=0;
   59803: out<=1;
   59804: out<=1;
   59805: out<=1;
   59806: out<=0;
   59807: out<=0;
   59808: out<=0;
   59809: out<=0;
   59810: out<=1;
   59811: out<=1;
   59812: out<=1;
   59813: out<=0;
   59814: out<=1;
   59815: out<=0;
   59816: out<=1;
   59817: out<=0;
   59818: out<=0;
   59819: out<=1;
   59820: out<=0;
   59821: out<=0;
   59822: out<=0;
   59823: out<=0;
   59824: out<=1;
   59825: out<=0;
   59826: out<=1;
   59827: out<=0;
   59828: out<=1;
   59829: out<=1;
   59830: out<=0;
   59831: out<=0;
   59832: out<=1;
   59833: out<=1;
   59834: out<=1;
   59835: out<=1;
   59836: out<=1;
   59837: out<=0;
   59838: out<=0;
   59839: out<=1;
   59840: out<=0;
   59841: out<=1;
   59842: out<=1;
   59843: out<=0;
   59844: out<=0;
   59845: out<=0;
   59846: out<=0;
   59847: out<=0;
   59848: out<=1;
   59849: out<=1;
   59850: out<=0;
   59851: out<=0;
   59852: out<=1;
   59853: out<=0;
   59854: out<=1;
   59855: out<=0;
   59856: out<=0;
   59857: out<=0;
   59858: out<=0;
   59859: out<=0;
   59860: out<=1;
   59861: out<=0;
   59862: out<=0;
   59863: out<=1;
   59864: out<=0;
   59865: out<=1;
   59866: out<=0;
   59867: out<=1;
   59868: out<=1;
   59869: out<=1;
   59870: out<=0;
   59871: out<=0;
   59872: out<=0;
   59873: out<=0;
   59874: out<=1;
   59875: out<=1;
   59876: out<=1;
   59877: out<=0;
   59878: out<=1;
   59879: out<=0;
   59880: out<=1;
   59881: out<=0;
   59882: out<=0;
   59883: out<=1;
   59884: out<=0;
   59885: out<=0;
   59886: out<=0;
   59887: out<=0;
   59888: out<=0;
   59889: out<=1;
   59890: out<=0;
   59891: out<=1;
   59892: out<=0;
   59893: out<=0;
   59894: out<=1;
   59895: out<=1;
   59896: out<=0;
   59897: out<=0;
   59898: out<=0;
   59899: out<=0;
   59900: out<=0;
   59901: out<=1;
   59902: out<=1;
   59903: out<=0;
   59904: out<=0;
   59905: out<=1;
   59906: out<=0;
   59907: out<=1;
   59908: out<=0;
   59909: out<=0;
   59910: out<=1;
   59911: out<=1;
   59912: out<=0;
   59913: out<=0;
   59914: out<=0;
   59915: out<=0;
   59916: out<=0;
   59917: out<=1;
   59918: out<=1;
   59919: out<=0;
   59920: out<=0;
   59921: out<=0;
   59922: out<=1;
   59923: out<=1;
   59924: out<=1;
   59925: out<=0;
   59926: out<=1;
   59927: out<=0;
   59928: out<=1;
   59929: out<=0;
   59930: out<=0;
   59931: out<=1;
   59932: out<=0;
   59933: out<=0;
   59934: out<=0;
   59935: out<=0;
   59936: out<=0;
   59937: out<=0;
   59938: out<=0;
   59939: out<=0;
   59940: out<=1;
   59941: out<=0;
   59942: out<=0;
   59943: out<=1;
   59944: out<=0;
   59945: out<=1;
   59946: out<=0;
   59947: out<=1;
   59948: out<=1;
   59949: out<=1;
   59950: out<=0;
   59951: out<=0;
   59952: out<=0;
   59953: out<=1;
   59954: out<=1;
   59955: out<=0;
   59956: out<=0;
   59957: out<=0;
   59958: out<=0;
   59959: out<=0;
   59960: out<=1;
   59961: out<=1;
   59962: out<=0;
   59963: out<=0;
   59964: out<=1;
   59965: out<=0;
   59966: out<=1;
   59967: out<=0;
   59968: out<=1;
   59969: out<=0;
   59970: out<=1;
   59971: out<=0;
   59972: out<=1;
   59973: out<=1;
   59974: out<=0;
   59975: out<=0;
   59976: out<=1;
   59977: out<=1;
   59978: out<=1;
   59979: out<=1;
   59980: out<=1;
   59981: out<=0;
   59982: out<=0;
   59983: out<=1;
   59984: out<=0;
   59985: out<=0;
   59986: out<=1;
   59987: out<=1;
   59988: out<=1;
   59989: out<=0;
   59990: out<=1;
   59991: out<=0;
   59992: out<=1;
   59993: out<=0;
   59994: out<=0;
   59995: out<=1;
   59996: out<=0;
   59997: out<=0;
   59998: out<=0;
   59999: out<=0;
   60000: out<=0;
   60001: out<=0;
   60002: out<=0;
   60003: out<=0;
   60004: out<=1;
   60005: out<=0;
   60006: out<=0;
   60007: out<=1;
   60008: out<=0;
   60009: out<=1;
   60010: out<=0;
   60011: out<=1;
   60012: out<=1;
   60013: out<=1;
   60014: out<=0;
   60015: out<=0;
   60016: out<=1;
   60017: out<=0;
   60018: out<=0;
   60019: out<=1;
   60020: out<=1;
   60021: out<=1;
   60022: out<=1;
   60023: out<=1;
   60024: out<=0;
   60025: out<=0;
   60026: out<=1;
   60027: out<=1;
   60028: out<=0;
   60029: out<=1;
   60030: out<=0;
   60031: out<=1;
   60032: out<=1;
   60033: out<=0;
   60034: out<=1;
   60035: out<=0;
   60036: out<=1;
   60037: out<=1;
   60038: out<=0;
   60039: out<=0;
   60040: out<=1;
   60041: out<=1;
   60042: out<=1;
   60043: out<=1;
   60044: out<=1;
   60045: out<=0;
   60046: out<=0;
   60047: out<=1;
   60048: out<=0;
   60049: out<=0;
   60050: out<=1;
   60051: out<=1;
   60052: out<=1;
   60053: out<=0;
   60054: out<=1;
   60055: out<=0;
   60056: out<=1;
   60057: out<=0;
   60058: out<=0;
   60059: out<=1;
   60060: out<=0;
   60061: out<=0;
   60062: out<=0;
   60063: out<=0;
   60064: out<=1;
   60065: out<=1;
   60066: out<=1;
   60067: out<=1;
   60068: out<=0;
   60069: out<=1;
   60070: out<=1;
   60071: out<=0;
   60072: out<=1;
   60073: out<=0;
   60074: out<=1;
   60075: out<=0;
   60076: out<=0;
   60077: out<=0;
   60078: out<=1;
   60079: out<=1;
   60080: out<=0;
   60081: out<=1;
   60082: out<=1;
   60083: out<=0;
   60084: out<=0;
   60085: out<=0;
   60086: out<=0;
   60087: out<=0;
   60088: out<=1;
   60089: out<=1;
   60090: out<=0;
   60091: out<=0;
   60092: out<=1;
   60093: out<=0;
   60094: out<=1;
   60095: out<=0;
   60096: out<=0;
   60097: out<=1;
   60098: out<=0;
   60099: out<=1;
   60100: out<=0;
   60101: out<=0;
   60102: out<=1;
   60103: out<=1;
   60104: out<=0;
   60105: out<=0;
   60106: out<=0;
   60107: out<=0;
   60108: out<=0;
   60109: out<=1;
   60110: out<=1;
   60111: out<=0;
   60112: out<=0;
   60113: out<=0;
   60114: out<=1;
   60115: out<=1;
   60116: out<=1;
   60117: out<=0;
   60118: out<=1;
   60119: out<=0;
   60120: out<=1;
   60121: out<=0;
   60122: out<=0;
   60123: out<=1;
   60124: out<=0;
   60125: out<=0;
   60126: out<=0;
   60127: out<=0;
   60128: out<=1;
   60129: out<=1;
   60130: out<=1;
   60131: out<=1;
   60132: out<=0;
   60133: out<=1;
   60134: out<=1;
   60135: out<=0;
   60136: out<=1;
   60137: out<=0;
   60138: out<=1;
   60139: out<=0;
   60140: out<=0;
   60141: out<=0;
   60142: out<=1;
   60143: out<=1;
   60144: out<=1;
   60145: out<=0;
   60146: out<=0;
   60147: out<=1;
   60148: out<=1;
   60149: out<=1;
   60150: out<=1;
   60151: out<=1;
   60152: out<=0;
   60153: out<=0;
   60154: out<=1;
   60155: out<=1;
   60156: out<=0;
   60157: out<=1;
   60158: out<=0;
   60159: out<=1;
   60160: out<=0;
   60161: out<=0;
   60162: out<=1;
   60163: out<=1;
   60164: out<=1;
   60165: out<=0;
   60166: out<=1;
   60167: out<=0;
   60168: out<=1;
   60169: out<=0;
   60170: out<=0;
   60171: out<=1;
   60172: out<=0;
   60173: out<=0;
   60174: out<=0;
   60175: out<=0;
   60176: out<=1;
   60177: out<=0;
   60178: out<=1;
   60179: out<=0;
   60180: out<=1;
   60181: out<=1;
   60182: out<=0;
   60183: out<=0;
   60184: out<=1;
   60185: out<=1;
   60186: out<=1;
   60187: out<=1;
   60188: out<=1;
   60189: out<=0;
   60190: out<=0;
   60191: out<=1;
   60192: out<=1;
   60193: out<=0;
   60194: out<=0;
   60195: out<=1;
   60196: out<=1;
   60197: out<=1;
   60198: out<=1;
   60199: out<=1;
   60200: out<=0;
   60201: out<=0;
   60202: out<=1;
   60203: out<=1;
   60204: out<=0;
   60205: out<=1;
   60206: out<=0;
   60207: out<=1;
   60208: out<=0;
   60209: out<=0;
   60210: out<=0;
   60211: out<=0;
   60212: out<=1;
   60213: out<=0;
   60214: out<=0;
   60215: out<=1;
   60216: out<=0;
   60217: out<=1;
   60218: out<=0;
   60219: out<=1;
   60220: out<=1;
   60221: out<=1;
   60222: out<=0;
   60223: out<=0;
   60224: out<=0;
   60225: out<=0;
   60226: out<=1;
   60227: out<=1;
   60228: out<=1;
   60229: out<=0;
   60230: out<=1;
   60231: out<=0;
   60232: out<=1;
   60233: out<=0;
   60234: out<=0;
   60235: out<=1;
   60236: out<=0;
   60237: out<=0;
   60238: out<=0;
   60239: out<=0;
   60240: out<=0;
   60241: out<=1;
   60242: out<=0;
   60243: out<=1;
   60244: out<=0;
   60245: out<=0;
   60246: out<=1;
   60247: out<=1;
   60248: out<=0;
   60249: out<=0;
   60250: out<=0;
   60251: out<=0;
   60252: out<=0;
   60253: out<=1;
   60254: out<=1;
   60255: out<=0;
   60256: out<=0;
   60257: out<=1;
   60258: out<=1;
   60259: out<=0;
   60260: out<=0;
   60261: out<=0;
   60262: out<=0;
   60263: out<=0;
   60264: out<=1;
   60265: out<=1;
   60266: out<=0;
   60267: out<=0;
   60268: out<=1;
   60269: out<=0;
   60270: out<=1;
   60271: out<=0;
   60272: out<=0;
   60273: out<=0;
   60274: out<=0;
   60275: out<=0;
   60276: out<=1;
   60277: out<=0;
   60278: out<=0;
   60279: out<=1;
   60280: out<=0;
   60281: out<=1;
   60282: out<=0;
   60283: out<=1;
   60284: out<=1;
   60285: out<=1;
   60286: out<=0;
   60287: out<=0;
   60288: out<=0;
   60289: out<=0;
   60290: out<=1;
   60291: out<=1;
   60292: out<=1;
   60293: out<=0;
   60294: out<=1;
   60295: out<=0;
   60296: out<=1;
   60297: out<=0;
   60298: out<=0;
   60299: out<=1;
   60300: out<=0;
   60301: out<=0;
   60302: out<=0;
   60303: out<=0;
   60304: out<=0;
   60305: out<=1;
   60306: out<=0;
   60307: out<=1;
   60308: out<=0;
   60309: out<=0;
   60310: out<=1;
   60311: out<=1;
   60312: out<=0;
   60313: out<=0;
   60314: out<=0;
   60315: out<=0;
   60316: out<=0;
   60317: out<=1;
   60318: out<=1;
   60319: out<=0;
   60320: out<=1;
   60321: out<=0;
   60322: out<=0;
   60323: out<=1;
   60324: out<=1;
   60325: out<=1;
   60326: out<=1;
   60327: out<=1;
   60328: out<=0;
   60329: out<=0;
   60330: out<=1;
   60331: out<=1;
   60332: out<=0;
   60333: out<=1;
   60334: out<=0;
   60335: out<=1;
   60336: out<=1;
   60337: out<=1;
   60338: out<=1;
   60339: out<=1;
   60340: out<=0;
   60341: out<=1;
   60342: out<=1;
   60343: out<=0;
   60344: out<=1;
   60345: out<=0;
   60346: out<=1;
   60347: out<=0;
   60348: out<=0;
   60349: out<=0;
   60350: out<=1;
   60351: out<=1;
   60352: out<=0;
   60353: out<=0;
   60354: out<=1;
   60355: out<=1;
   60356: out<=1;
   60357: out<=0;
   60358: out<=1;
   60359: out<=0;
   60360: out<=1;
   60361: out<=0;
   60362: out<=0;
   60363: out<=1;
   60364: out<=0;
   60365: out<=0;
   60366: out<=0;
   60367: out<=0;
   60368: out<=1;
   60369: out<=0;
   60370: out<=1;
   60371: out<=0;
   60372: out<=1;
   60373: out<=1;
   60374: out<=0;
   60375: out<=0;
   60376: out<=1;
   60377: out<=1;
   60378: out<=1;
   60379: out<=1;
   60380: out<=1;
   60381: out<=0;
   60382: out<=0;
   60383: out<=1;
   60384: out<=0;
   60385: out<=1;
   60386: out<=1;
   60387: out<=0;
   60388: out<=0;
   60389: out<=0;
   60390: out<=0;
   60391: out<=0;
   60392: out<=1;
   60393: out<=1;
   60394: out<=0;
   60395: out<=0;
   60396: out<=1;
   60397: out<=0;
   60398: out<=1;
   60399: out<=0;
   60400: out<=1;
   60401: out<=1;
   60402: out<=1;
   60403: out<=1;
   60404: out<=0;
   60405: out<=1;
   60406: out<=1;
   60407: out<=0;
   60408: out<=1;
   60409: out<=0;
   60410: out<=1;
   60411: out<=0;
   60412: out<=0;
   60413: out<=0;
   60414: out<=1;
   60415: out<=1;
   60416: out<=0;
   60417: out<=1;
   60418: out<=1;
   60419: out<=0;
   60420: out<=1;
   60421: out<=1;
   60422: out<=1;
   60423: out<=1;
   60424: out<=0;
   60425: out<=0;
   60426: out<=1;
   60427: out<=1;
   60428: out<=1;
   60429: out<=0;
   60430: out<=1;
   60431: out<=0;
   60432: out<=1;
   60433: out<=1;
   60434: out<=1;
   60435: out<=1;
   60436: out<=1;
   60437: out<=0;
   60438: out<=0;
   60439: out<=1;
   60440: out<=0;
   60441: out<=1;
   60442: out<=0;
   60443: out<=1;
   60444: out<=0;
   60445: out<=0;
   60446: out<=1;
   60447: out<=1;
   60448: out<=0;
   60449: out<=0;
   60450: out<=1;
   60451: out<=1;
   60452: out<=0;
   60453: out<=1;
   60454: out<=0;
   60455: out<=1;
   60456: out<=0;
   60457: out<=1;
   60458: out<=1;
   60459: out<=0;
   60460: out<=0;
   60461: out<=0;
   60462: out<=0;
   60463: out<=0;
   60464: out<=1;
   60465: out<=0;
   60466: out<=1;
   60467: out<=0;
   60468: out<=0;
   60469: out<=0;
   60470: out<=1;
   60471: out<=1;
   60472: out<=0;
   60473: out<=0;
   60474: out<=0;
   60475: out<=0;
   60476: out<=1;
   60477: out<=0;
   60478: out<=0;
   60479: out<=1;
   60480: out<=1;
   60481: out<=0;
   60482: out<=0;
   60483: out<=1;
   60484: out<=0;
   60485: out<=0;
   60486: out<=0;
   60487: out<=0;
   60488: out<=1;
   60489: out<=1;
   60490: out<=0;
   60491: out<=0;
   60492: out<=0;
   60493: out<=1;
   60494: out<=0;
   60495: out<=1;
   60496: out<=1;
   60497: out<=1;
   60498: out<=1;
   60499: out<=1;
   60500: out<=1;
   60501: out<=0;
   60502: out<=0;
   60503: out<=1;
   60504: out<=0;
   60505: out<=1;
   60506: out<=0;
   60507: out<=1;
   60508: out<=0;
   60509: out<=0;
   60510: out<=1;
   60511: out<=1;
   60512: out<=0;
   60513: out<=0;
   60514: out<=1;
   60515: out<=1;
   60516: out<=0;
   60517: out<=1;
   60518: out<=0;
   60519: out<=1;
   60520: out<=0;
   60521: out<=1;
   60522: out<=1;
   60523: out<=0;
   60524: out<=0;
   60525: out<=0;
   60526: out<=0;
   60527: out<=0;
   60528: out<=0;
   60529: out<=1;
   60530: out<=0;
   60531: out<=1;
   60532: out<=1;
   60533: out<=1;
   60534: out<=0;
   60535: out<=0;
   60536: out<=1;
   60537: out<=1;
   60538: out<=1;
   60539: out<=1;
   60540: out<=0;
   60541: out<=1;
   60542: out<=1;
   60543: out<=0;
   60544: out<=0;
   60545: out<=1;
   60546: out<=1;
   60547: out<=0;
   60548: out<=1;
   60549: out<=1;
   60550: out<=1;
   60551: out<=1;
   60552: out<=0;
   60553: out<=0;
   60554: out<=1;
   60555: out<=1;
   60556: out<=1;
   60557: out<=0;
   60558: out<=1;
   60559: out<=0;
   60560: out<=0;
   60561: out<=0;
   60562: out<=0;
   60563: out<=0;
   60564: out<=0;
   60565: out<=1;
   60566: out<=1;
   60567: out<=0;
   60568: out<=1;
   60569: out<=0;
   60570: out<=1;
   60571: out<=0;
   60572: out<=1;
   60573: out<=1;
   60574: out<=0;
   60575: out<=0;
   60576: out<=0;
   60577: out<=0;
   60578: out<=1;
   60579: out<=1;
   60580: out<=0;
   60581: out<=1;
   60582: out<=0;
   60583: out<=1;
   60584: out<=0;
   60585: out<=1;
   60586: out<=1;
   60587: out<=0;
   60588: out<=0;
   60589: out<=0;
   60590: out<=0;
   60591: out<=0;
   60592: out<=0;
   60593: out<=1;
   60594: out<=0;
   60595: out<=1;
   60596: out<=1;
   60597: out<=1;
   60598: out<=0;
   60599: out<=0;
   60600: out<=1;
   60601: out<=1;
   60602: out<=1;
   60603: out<=1;
   60604: out<=0;
   60605: out<=1;
   60606: out<=1;
   60607: out<=0;
   60608: out<=1;
   60609: out<=0;
   60610: out<=0;
   60611: out<=1;
   60612: out<=0;
   60613: out<=0;
   60614: out<=0;
   60615: out<=0;
   60616: out<=1;
   60617: out<=1;
   60618: out<=0;
   60619: out<=0;
   60620: out<=0;
   60621: out<=1;
   60622: out<=0;
   60623: out<=1;
   60624: out<=0;
   60625: out<=0;
   60626: out<=0;
   60627: out<=0;
   60628: out<=0;
   60629: out<=1;
   60630: out<=1;
   60631: out<=0;
   60632: out<=1;
   60633: out<=0;
   60634: out<=1;
   60635: out<=0;
   60636: out<=1;
   60637: out<=1;
   60638: out<=0;
   60639: out<=0;
   60640: out<=0;
   60641: out<=0;
   60642: out<=1;
   60643: out<=1;
   60644: out<=0;
   60645: out<=1;
   60646: out<=0;
   60647: out<=1;
   60648: out<=0;
   60649: out<=1;
   60650: out<=1;
   60651: out<=0;
   60652: out<=0;
   60653: out<=0;
   60654: out<=0;
   60655: out<=0;
   60656: out<=1;
   60657: out<=0;
   60658: out<=1;
   60659: out<=0;
   60660: out<=0;
   60661: out<=0;
   60662: out<=1;
   60663: out<=1;
   60664: out<=0;
   60665: out<=0;
   60666: out<=0;
   60667: out<=0;
   60668: out<=1;
   60669: out<=0;
   60670: out<=0;
   60671: out<=1;
   60672: out<=1;
   60673: out<=1;
   60674: out<=1;
   60675: out<=1;
   60676: out<=1;
   60677: out<=0;
   60678: out<=0;
   60679: out<=1;
   60680: out<=0;
   60681: out<=1;
   60682: out<=0;
   60683: out<=1;
   60684: out<=0;
   60685: out<=0;
   60686: out<=1;
   60687: out<=1;
   60688: out<=1;
   60689: out<=0;
   60690: out<=0;
   60691: out<=1;
   60692: out<=0;
   60693: out<=0;
   60694: out<=0;
   60695: out<=0;
   60696: out<=1;
   60697: out<=1;
   60698: out<=0;
   60699: out<=0;
   60700: out<=0;
   60701: out<=1;
   60702: out<=0;
   60703: out<=1;
   60704: out<=0;
   60705: out<=1;
   60706: out<=0;
   60707: out<=1;
   60708: out<=1;
   60709: out<=1;
   60710: out<=0;
   60711: out<=0;
   60712: out<=1;
   60713: out<=1;
   60714: out<=1;
   60715: out<=1;
   60716: out<=0;
   60717: out<=1;
   60718: out<=1;
   60719: out<=0;
   60720: out<=0;
   60721: out<=0;
   60722: out<=1;
   60723: out<=1;
   60724: out<=0;
   60725: out<=1;
   60726: out<=0;
   60727: out<=1;
   60728: out<=0;
   60729: out<=1;
   60730: out<=1;
   60731: out<=0;
   60732: out<=0;
   60733: out<=0;
   60734: out<=0;
   60735: out<=0;
   60736: out<=1;
   60737: out<=1;
   60738: out<=1;
   60739: out<=1;
   60740: out<=1;
   60741: out<=0;
   60742: out<=0;
   60743: out<=1;
   60744: out<=0;
   60745: out<=1;
   60746: out<=0;
   60747: out<=1;
   60748: out<=0;
   60749: out<=0;
   60750: out<=1;
   60751: out<=1;
   60752: out<=0;
   60753: out<=1;
   60754: out<=1;
   60755: out<=0;
   60756: out<=1;
   60757: out<=1;
   60758: out<=1;
   60759: out<=1;
   60760: out<=0;
   60761: out<=0;
   60762: out<=1;
   60763: out<=1;
   60764: out<=1;
   60765: out<=0;
   60766: out<=1;
   60767: out<=0;
   60768: out<=1;
   60769: out<=0;
   60770: out<=1;
   60771: out<=0;
   60772: out<=0;
   60773: out<=0;
   60774: out<=1;
   60775: out<=1;
   60776: out<=0;
   60777: out<=0;
   60778: out<=0;
   60779: out<=0;
   60780: out<=1;
   60781: out<=0;
   60782: out<=0;
   60783: out<=1;
   60784: out<=0;
   60785: out<=0;
   60786: out<=1;
   60787: out<=1;
   60788: out<=0;
   60789: out<=1;
   60790: out<=0;
   60791: out<=1;
   60792: out<=0;
   60793: out<=1;
   60794: out<=1;
   60795: out<=0;
   60796: out<=0;
   60797: out<=0;
   60798: out<=0;
   60799: out<=0;
   60800: out<=0;
   60801: out<=0;
   60802: out<=0;
   60803: out<=0;
   60804: out<=0;
   60805: out<=1;
   60806: out<=1;
   60807: out<=0;
   60808: out<=1;
   60809: out<=0;
   60810: out<=1;
   60811: out<=0;
   60812: out<=1;
   60813: out<=1;
   60814: out<=0;
   60815: out<=0;
   60816: out<=1;
   60817: out<=0;
   60818: out<=0;
   60819: out<=1;
   60820: out<=0;
   60821: out<=0;
   60822: out<=0;
   60823: out<=0;
   60824: out<=1;
   60825: out<=1;
   60826: out<=0;
   60827: out<=0;
   60828: out<=0;
   60829: out<=1;
   60830: out<=0;
   60831: out<=1;
   60832: out<=1;
   60833: out<=0;
   60834: out<=1;
   60835: out<=0;
   60836: out<=0;
   60837: out<=0;
   60838: out<=1;
   60839: out<=1;
   60840: out<=0;
   60841: out<=0;
   60842: out<=0;
   60843: out<=0;
   60844: out<=1;
   60845: out<=0;
   60846: out<=0;
   60847: out<=1;
   60848: out<=0;
   60849: out<=0;
   60850: out<=1;
   60851: out<=1;
   60852: out<=0;
   60853: out<=1;
   60854: out<=0;
   60855: out<=1;
   60856: out<=0;
   60857: out<=1;
   60858: out<=1;
   60859: out<=0;
   60860: out<=0;
   60861: out<=0;
   60862: out<=0;
   60863: out<=0;
   60864: out<=0;
   60865: out<=0;
   60866: out<=0;
   60867: out<=0;
   60868: out<=0;
   60869: out<=1;
   60870: out<=1;
   60871: out<=0;
   60872: out<=1;
   60873: out<=0;
   60874: out<=1;
   60875: out<=0;
   60876: out<=1;
   60877: out<=1;
   60878: out<=0;
   60879: out<=0;
   60880: out<=0;
   60881: out<=1;
   60882: out<=1;
   60883: out<=0;
   60884: out<=1;
   60885: out<=1;
   60886: out<=1;
   60887: out<=1;
   60888: out<=0;
   60889: out<=0;
   60890: out<=1;
   60891: out<=1;
   60892: out<=1;
   60893: out<=0;
   60894: out<=1;
   60895: out<=0;
   60896: out<=0;
   60897: out<=1;
   60898: out<=0;
   60899: out<=1;
   60900: out<=1;
   60901: out<=1;
   60902: out<=0;
   60903: out<=0;
   60904: out<=1;
   60905: out<=1;
   60906: out<=1;
   60907: out<=1;
   60908: out<=0;
   60909: out<=1;
   60910: out<=1;
   60911: out<=0;
   60912: out<=0;
   60913: out<=0;
   60914: out<=1;
   60915: out<=1;
   60916: out<=0;
   60917: out<=1;
   60918: out<=0;
   60919: out<=1;
   60920: out<=0;
   60921: out<=1;
   60922: out<=1;
   60923: out<=0;
   60924: out<=0;
   60925: out<=0;
   60926: out<=0;
   60927: out<=0;
   60928: out<=0;
   60929: out<=0;
   60930: out<=1;
   60931: out<=1;
   60932: out<=0;
   60933: out<=1;
   60934: out<=0;
   60935: out<=1;
   60936: out<=0;
   60937: out<=1;
   60938: out<=1;
   60939: out<=0;
   60940: out<=0;
   60941: out<=0;
   60942: out<=0;
   60943: out<=0;
   60944: out<=0;
   60945: out<=1;
   60946: out<=0;
   60947: out<=1;
   60948: out<=1;
   60949: out<=1;
   60950: out<=0;
   60951: out<=0;
   60952: out<=1;
   60953: out<=1;
   60954: out<=1;
   60955: out<=1;
   60956: out<=0;
   60957: out<=1;
   60958: out<=1;
   60959: out<=0;
   60960: out<=0;
   60961: out<=1;
   60962: out<=1;
   60963: out<=0;
   60964: out<=1;
   60965: out<=1;
   60966: out<=1;
   60967: out<=1;
   60968: out<=0;
   60969: out<=0;
   60970: out<=1;
   60971: out<=1;
   60972: out<=1;
   60973: out<=0;
   60974: out<=1;
   60975: out<=0;
   60976: out<=0;
   60977: out<=0;
   60978: out<=0;
   60979: out<=0;
   60980: out<=0;
   60981: out<=1;
   60982: out<=1;
   60983: out<=0;
   60984: out<=1;
   60985: out<=0;
   60986: out<=1;
   60987: out<=0;
   60988: out<=1;
   60989: out<=1;
   60990: out<=0;
   60991: out<=0;
   60992: out<=0;
   60993: out<=0;
   60994: out<=1;
   60995: out<=1;
   60996: out<=0;
   60997: out<=1;
   60998: out<=0;
   60999: out<=1;
   61000: out<=0;
   61001: out<=1;
   61002: out<=1;
   61003: out<=0;
   61004: out<=0;
   61005: out<=0;
   61006: out<=0;
   61007: out<=0;
   61008: out<=1;
   61009: out<=0;
   61010: out<=1;
   61011: out<=0;
   61012: out<=0;
   61013: out<=0;
   61014: out<=1;
   61015: out<=1;
   61016: out<=0;
   61017: out<=0;
   61018: out<=0;
   61019: out<=0;
   61020: out<=1;
   61021: out<=0;
   61022: out<=0;
   61023: out<=1;
   61024: out<=1;
   61025: out<=0;
   61026: out<=0;
   61027: out<=1;
   61028: out<=0;
   61029: out<=0;
   61030: out<=0;
   61031: out<=0;
   61032: out<=1;
   61033: out<=1;
   61034: out<=0;
   61035: out<=0;
   61036: out<=0;
   61037: out<=1;
   61038: out<=0;
   61039: out<=1;
   61040: out<=0;
   61041: out<=0;
   61042: out<=0;
   61043: out<=0;
   61044: out<=0;
   61045: out<=1;
   61046: out<=1;
   61047: out<=0;
   61048: out<=1;
   61049: out<=0;
   61050: out<=1;
   61051: out<=0;
   61052: out<=1;
   61053: out<=1;
   61054: out<=0;
   61055: out<=0;
   61056: out<=0;
   61057: out<=0;
   61058: out<=1;
   61059: out<=1;
   61060: out<=0;
   61061: out<=1;
   61062: out<=0;
   61063: out<=1;
   61064: out<=0;
   61065: out<=1;
   61066: out<=1;
   61067: out<=0;
   61068: out<=0;
   61069: out<=0;
   61070: out<=0;
   61071: out<=0;
   61072: out<=1;
   61073: out<=0;
   61074: out<=1;
   61075: out<=0;
   61076: out<=0;
   61077: out<=0;
   61078: out<=1;
   61079: out<=1;
   61080: out<=0;
   61081: out<=0;
   61082: out<=0;
   61083: out<=0;
   61084: out<=1;
   61085: out<=0;
   61086: out<=0;
   61087: out<=1;
   61088: out<=0;
   61089: out<=1;
   61090: out<=1;
   61091: out<=0;
   61092: out<=1;
   61093: out<=1;
   61094: out<=1;
   61095: out<=1;
   61096: out<=0;
   61097: out<=0;
   61098: out<=1;
   61099: out<=1;
   61100: out<=1;
   61101: out<=0;
   61102: out<=1;
   61103: out<=0;
   61104: out<=1;
   61105: out<=1;
   61106: out<=1;
   61107: out<=1;
   61108: out<=1;
   61109: out<=0;
   61110: out<=0;
   61111: out<=1;
   61112: out<=0;
   61113: out<=1;
   61114: out<=0;
   61115: out<=1;
   61116: out<=0;
   61117: out<=0;
   61118: out<=1;
   61119: out<=1;
   61120: out<=0;
   61121: out<=0;
   61122: out<=1;
   61123: out<=1;
   61124: out<=0;
   61125: out<=1;
   61126: out<=0;
   61127: out<=1;
   61128: out<=0;
   61129: out<=1;
   61130: out<=1;
   61131: out<=0;
   61132: out<=0;
   61133: out<=0;
   61134: out<=0;
   61135: out<=0;
   61136: out<=0;
   61137: out<=1;
   61138: out<=0;
   61139: out<=1;
   61140: out<=1;
   61141: out<=1;
   61142: out<=0;
   61143: out<=0;
   61144: out<=1;
   61145: out<=1;
   61146: out<=1;
   61147: out<=1;
   61148: out<=0;
   61149: out<=1;
   61150: out<=1;
   61151: out<=0;
   61152: out<=1;
   61153: out<=0;
   61154: out<=0;
   61155: out<=1;
   61156: out<=0;
   61157: out<=0;
   61158: out<=0;
   61159: out<=0;
   61160: out<=1;
   61161: out<=1;
   61162: out<=0;
   61163: out<=0;
   61164: out<=0;
   61165: out<=1;
   61166: out<=0;
   61167: out<=1;
   61168: out<=1;
   61169: out<=1;
   61170: out<=1;
   61171: out<=1;
   61172: out<=1;
   61173: out<=0;
   61174: out<=0;
   61175: out<=1;
   61176: out<=0;
   61177: out<=1;
   61178: out<=0;
   61179: out<=1;
   61180: out<=0;
   61181: out<=0;
   61182: out<=1;
   61183: out<=1;
   61184: out<=1;
   61185: out<=0;
   61186: out<=1;
   61187: out<=0;
   61188: out<=0;
   61189: out<=0;
   61190: out<=1;
   61191: out<=1;
   61192: out<=0;
   61193: out<=0;
   61194: out<=0;
   61195: out<=0;
   61196: out<=1;
   61197: out<=0;
   61198: out<=0;
   61199: out<=1;
   61200: out<=0;
   61201: out<=0;
   61202: out<=1;
   61203: out<=1;
   61204: out<=0;
   61205: out<=1;
   61206: out<=0;
   61207: out<=1;
   61208: out<=0;
   61209: out<=1;
   61210: out<=1;
   61211: out<=0;
   61212: out<=0;
   61213: out<=0;
   61214: out<=0;
   61215: out<=0;
   61216: out<=0;
   61217: out<=0;
   61218: out<=0;
   61219: out<=0;
   61220: out<=0;
   61221: out<=1;
   61222: out<=1;
   61223: out<=0;
   61224: out<=1;
   61225: out<=0;
   61226: out<=1;
   61227: out<=0;
   61228: out<=1;
   61229: out<=1;
   61230: out<=0;
   61231: out<=0;
   61232: out<=1;
   61233: out<=0;
   61234: out<=0;
   61235: out<=1;
   61236: out<=0;
   61237: out<=0;
   61238: out<=0;
   61239: out<=0;
   61240: out<=1;
   61241: out<=1;
   61242: out<=0;
   61243: out<=0;
   61244: out<=0;
   61245: out<=1;
   61246: out<=0;
   61247: out<=1;
   61248: out<=0;
   61249: out<=1;
   61250: out<=0;
   61251: out<=1;
   61252: out<=1;
   61253: out<=1;
   61254: out<=0;
   61255: out<=0;
   61256: out<=1;
   61257: out<=1;
   61258: out<=1;
   61259: out<=1;
   61260: out<=0;
   61261: out<=1;
   61262: out<=1;
   61263: out<=0;
   61264: out<=0;
   61265: out<=0;
   61266: out<=1;
   61267: out<=1;
   61268: out<=0;
   61269: out<=1;
   61270: out<=0;
   61271: out<=1;
   61272: out<=0;
   61273: out<=1;
   61274: out<=1;
   61275: out<=0;
   61276: out<=0;
   61277: out<=0;
   61278: out<=0;
   61279: out<=0;
   61280: out<=0;
   61281: out<=0;
   61282: out<=0;
   61283: out<=0;
   61284: out<=0;
   61285: out<=1;
   61286: out<=1;
   61287: out<=0;
   61288: out<=1;
   61289: out<=0;
   61290: out<=1;
   61291: out<=0;
   61292: out<=1;
   61293: out<=1;
   61294: out<=0;
   61295: out<=0;
   61296: out<=0;
   61297: out<=1;
   61298: out<=1;
   61299: out<=0;
   61300: out<=1;
   61301: out<=1;
   61302: out<=1;
   61303: out<=1;
   61304: out<=0;
   61305: out<=0;
   61306: out<=1;
   61307: out<=1;
   61308: out<=1;
   61309: out<=0;
   61310: out<=1;
   61311: out<=0;
   61312: out<=0;
   61313: out<=1;
   61314: out<=0;
   61315: out<=1;
   61316: out<=1;
   61317: out<=1;
   61318: out<=0;
   61319: out<=0;
   61320: out<=1;
   61321: out<=1;
   61322: out<=1;
   61323: out<=1;
   61324: out<=0;
   61325: out<=1;
   61326: out<=1;
   61327: out<=0;
   61328: out<=0;
   61329: out<=0;
   61330: out<=1;
   61331: out<=1;
   61332: out<=0;
   61333: out<=1;
   61334: out<=0;
   61335: out<=1;
   61336: out<=0;
   61337: out<=1;
   61338: out<=1;
   61339: out<=0;
   61340: out<=0;
   61341: out<=0;
   61342: out<=0;
   61343: out<=0;
   61344: out<=1;
   61345: out<=1;
   61346: out<=1;
   61347: out<=1;
   61348: out<=1;
   61349: out<=0;
   61350: out<=0;
   61351: out<=1;
   61352: out<=0;
   61353: out<=1;
   61354: out<=0;
   61355: out<=1;
   61356: out<=0;
   61357: out<=0;
   61358: out<=1;
   61359: out<=1;
   61360: out<=1;
   61361: out<=0;
   61362: out<=0;
   61363: out<=1;
   61364: out<=0;
   61365: out<=0;
   61366: out<=0;
   61367: out<=0;
   61368: out<=1;
   61369: out<=1;
   61370: out<=0;
   61371: out<=0;
   61372: out<=0;
   61373: out<=1;
   61374: out<=0;
   61375: out<=1;
   61376: out<=1;
   61377: out<=0;
   61378: out<=1;
   61379: out<=0;
   61380: out<=0;
   61381: out<=0;
   61382: out<=1;
   61383: out<=1;
   61384: out<=0;
   61385: out<=0;
   61386: out<=0;
   61387: out<=0;
   61388: out<=1;
   61389: out<=0;
   61390: out<=0;
   61391: out<=1;
   61392: out<=0;
   61393: out<=0;
   61394: out<=1;
   61395: out<=1;
   61396: out<=0;
   61397: out<=1;
   61398: out<=0;
   61399: out<=1;
   61400: out<=0;
   61401: out<=1;
   61402: out<=1;
   61403: out<=0;
   61404: out<=0;
   61405: out<=0;
   61406: out<=0;
   61407: out<=0;
   61408: out<=1;
   61409: out<=1;
   61410: out<=1;
   61411: out<=1;
   61412: out<=1;
   61413: out<=0;
   61414: out<=0;
   61415: out<=1;
   61416: out<=0;
   61417: out<=1;
   61418: out<=0;
   61419: out<=1;
   61420: out<=0;
   61421: out<=0;
   61422: out<=1;
   61423: out<=1;
   61424: out<=0;
   61425: out<=1;
   61426: out<=1;
   61427: out<=0;
   61428: out<=1;
   61429: out<=1;
   61430: out<=1;
   61431: out<=1;
   61432: out<=0;
   61433: out<=0;
   61434: out<=1;
   61435: out<=1;
   61436: out<=1;
   61437: out<=0;
   61438: out<=1;
   61439: out<=0;
   61440: out<=1;
   61441: out<=0;
   61442: out<=1;
   61443: out<=0;
   61444: out<=1;
   61445: out<=1;
   61446: out<=0;
   61447: out<=0;
   61448: out<=0;
   61449: out<=0;
   61450: out<=0;
   61451: out<=0;
   61452: out<=0;
   61453: out<=1;
   61454: out<=1;
   61455: out<=0;
   61456: out<=0;
   61457: out<=0;
   61458: out<=1;
   61459: out<=1;
   61460: out<=1;
   61461: out<=0;
   61462: out<=1;
   61463: out<=0;
   61464: out<=0;
   61465: out<=1;
   61466: out<=1;
   61467: out<=0;
   61468: out<=1;
   61469: out<=1;
   61470: out<=1;
   61471: out<=1;
   61472: out<=1;
   61473: out<=1;
   61474: out<=1;
   61475: out<=1;
   61476: out<=0;
   61477: out<=1;
   61478: out<=1;
   61479: out<=0;
   61480: out<=0;
   61481: out<=1;
   61482: out<=0;
   61483: out<=1;
   61484: out<=1;
   61485: out<=1;
   61486: out<=0;
   61487: out<=0;
   61488: out<=0;
   61489: out<=1;
   61490: out<=1;
   61491: out<=0;
   61492: out<=0;
   61493: out<=0;
   61494: out<=0;
   61495: out<=0;
   61496: out<=0;
   61497: out<=0;
   61498: out<=1;
   61499: out<=1;
   61500: out<=0;
   61501: out<=1;
   61502: out<=0;
   61503: out<=1;
   61504: out<=0;
   61505: out<=1;
   61506: out<=0;
   61507: out<=1;
   61508: out<=0;
   61509: out<=0;
   61510: out<=1;
   61511: out<=1;
   61512: out<=1;
   61513: out<=1;
   61514: out<=1;
   61515: out<=1;
   61516: out<=1;
   61517: out<=0;
   61518: out<=0;
   61519: out<=1;
   61520: out<=0;
   61521: out<=0;
   61522: out<=1;
   61523: out<=1;
   61524: out<=1;
   61525: out<=0;
   61526: out<=1;
   61527: out<=0;
   61528: out<=0;
   61529: out<=1;
   61530: out<=1;
   61531: out<=0;
   61532: out<=1;
   61533: out<=1;
   61534: out<=1;
   61535: out<=1;
   61536: out<=1;
   61537: out<=1;
   61538: out<=1;
   61539: out<=1;
   61540: out<=0;
   61541: out<=1;
   61542: out<=1;
   61543: out<=0;
   61544: out<=0;
   61545: out<=1;
   61546: out<=0;
   61547: out<=1;
   61548: out<=1;
   61549: out<=1;
   61550: out<=0;
   61551: out<=0;
   61552: out<=1;
   61553: out<=0;
   61554: out<=0;
   61555: out<=1;
   61556: out<=1;
   61557: out<=1;
   61558: out<=1;
   61559: out<=1;
   61560: out<=1;
   61561: out<=1;
   61562: out<=0;
   61563: out<=0;
   61564: out<=1;
   61565: out<=0;
   61566: out<=1;
   61567: out<=0;
   61568: out<=0;
   61569: out<=1;
   61570: out<=0;
   61571: out<=1;
   61572: out<=0;
   61573: out<=0;
   61574: out<=1;
   61575: out<=1;
   61576: out<=1;
   61577: out<=1;
   61578: out<=1;
   61579: out<=1;
   61580: out<=1;
   61581: out<=0;
   61582: out<=0;
   61583: out<=1;
   61584: out<=0;
   61585: out<=0;
   61586: out<=1;
   61587: out<=1;
   61588: out<=1;
   61589: out<=0;
   61590: out<=1;
   61591: out<=0;
   61592: out<=0;
   61593: out<=1;
   61594: out<=1;
   61595: out<=0;
   61596: out<=1;
   61597: out<=1;
   61598: out<=1;
   61599: out<=1;
   61600: out<=0;
   61601: out<=0;
   61602: out<=0;
   61603: out<=0;
   61604: out<=1;
   61605: out<=0;
   61606: out<=0;
   61607: out<=1;
   61608: out<=1;
   61609: out<=0;
   61610: out<=1;
   61611: out<=0;
   61612: out<=0;
   61613: out<=0;
   61614: out<=1;
   61615: out<=1;
   61616: out<=0;
   61617: out<=1;
   61618: out<=1;
   61619: out<=0;
   61620: out<=0;
   61621: out<=0;
   61622: out<=0;
   61623: out<=0;
   61624: out<=0;
   61625: out<=0;
   61626: out<=1;
   61627: out<=1;
   61628: out<=0;
   61629: out<=1;
   61630: out<=0;
   61631: out<=1;
   61632: out<=1;
   61633: out<=0;
   61634: out<=1;
   61635: out<=0;
   61636: out<=1;
   61637: out<=1;
   61638: out<=0;
   61639: out<=0;
   61640: out<=0;
   61641: out<=0;
   61642: out<=0;
   61643: out<=0;
   61644: out<=0;
   61645: out<=1;
   61646: out<=1;
   61647: out<=0;
   61648: out<=0;
   61649: out<=0;
   61650: out<=1;
   61651: out<=1;
   61652: out<=1;
   61653: out<=0;
   61654: out<=1;
   61655: out<=0;
   61656: out<=0;
   61657: out<=1;
   61658: out<=1;
   61659: out<=0;
   61660: out<=1;
   61661: out<=1;
   61662: out<=1;
   61663: out<=1;
   61664: out<=0;
   61665: out<=0;
   61666: out<=0;
   61667: out<=0;
   61668: out<=1;
   61669: out<=0;
   61670: out<=0;
   61671: out<=1;
   61672: out<=1;
   61673: out<=0;
   61674: out<=1;
   61675: out<=0;
   61676: out<=0;
   61677: out<=0;
   61678: out<=1;
   61679: out<=1;
   61680: out<=1;
   61681: out<=0;
   61682: out<=0;
   61683: out<=1;
   61684: out<=1;
   61685: out<=1;
   61686: out<=1;
   61687: out<=1;
   61688: out<=1;
   61689: out<=1;
   61690: out<=0;
   61691: out<=0;
   61692: out<=1;
   61693: out<=0;
   61694: out<=1;
   61695: out<=0;
   61696: out<=0;
   61697: out<=0;
   61698: out<=1;
   61699: out<=1;
   61700: out<=1;
   61701: out<=0;
   61702: out<=1;
   61703: out<=0;
   61704: out<=0;
   61705: out<=1;
   61706: out<=1;
   61707: out<=0;
   61708: out<=1;
   61709: out<=1;
   61710: out<=1;
   61711: out<=1;
   61712: out<=0;
   61713: out<=1;
   61714: out<=0;
   61715: out<=1;
   61716: out<=0;
   61717: out<=0;
   61718: out<=1;
   61719: out<=1;
   61720: out<=1;
   61721: out<=1;
   61722: out<=1;
   61723: out<=1;
   61724: out<=1;
   61725: out<=0;
   61726: out<=0;
   61727: out<=1;
   61728: out<=1;
   61729: out<=0;
   61730: out<=0;
   61731: out<=1;
   61732: out<=1;
   61733: out<=1;
   61734: out<=1;
   61735: out<=1;
   61736: out<=1;
   61737: out<=1;
   61738: out<=0;
   61739: out<=0;
   61740: out<=1;
   61741: out<=0;
   61742: out<=1;
   61743: out<=0;
   61744: out<=1;
   61745: out<=1;
   61746: out<=1;
   61747: out<=1;
   61748: out<=0;
   61749: out<=1;
   61750: out<=1;
   61751: out<=0;
   61752: out<=0;
   61753: out<=1;
   61754: out<=0;
   61755: out<=1;
   61756: out<=1;
   61757: out<=1;
   61758: out<=0;
   61759: out<=0;
   61760: out<=0;
   61761: out<=0;
   61762: out<=1;
   61763: out<=1;
   61764: out<=1;
   61765: out<=0;
   61766: out<=1;
   61767: out<=0;
   61768: out<=0;
   61769: out<=1;
   61770: out<=1;
   61771: out<=0;
   61772: out<=1;
   61773: out<=1;
   61774: out<=1;
   61775: out<=1;
   61776: out<=1;
   61777: out<=0;
   61778: out<=1;
   61779: out<=0;
   61780: out<=1;
   61781: out<=1;
   61782: out<=0;
   61783: out<=0;
   61784: out<=0;
   61785: out<=0;
   61786: out<=0;
   61787: out<=0;
   61788: out<=0;
   61789: out<=1;
   61790: out<=1;
   61791: out<=0;
   61792: out<=0;
   61793: out<=1;
   61794: out<=1;
   61795: out<=0;
   61796: out<=0;
   61797: out<=0;
   61798: out<=0;
   61799: out<=0;
   61800: out<=0;
   61801: out<=0;
   61802: out<=1;
   61803: out<=1;
   61804: out<=0;
   61805: out<=1;
   61806: out<=0;
   61807: out<=1;
   61808: out<=1;
   61809: out<=1;
   61810: out<=1;
   61811: out<=1;
   61812: out<=0;
   61813: out<=1;
   61814: out<=1;
   61815: out<=0;
   61816: out<=0;
   61817: out<=1;
   61818: out<=0;
   61819: out<=1;
   61820: out<=1;
   61821: out<=1;
   61822: out<=0;
   61823: out<=0;
   61824: out<=0;
   61825: out<=0;
   61826: out<=1;
   61827: out<=1;
   61828: out<=1;
   61829: out<=0;
   61830: out<=1;
   61831: out<=0;
   61832: out<=0;
   61833: out<=1;
   61834: out<=1;
   61835: out<=0;
   61836: out<=1;
   61837: out<=1;
   61838: out<=1;
   61839: out<=1;
   61840: out<=1;
   61841: out<=0;
   61842: out<=1;
   61843: out<=0;
   61844: out<=1;
   61845: out<=1;
   61846: out<=0;
   61847: out<=0;
   61848: out<=0;
   61849: out<=0;
   61850: out<=0;
   61851: out<=0;
   61852: out<=0;
   61853: out<=1;
   61854: out<=1;
   61855: out<=0;
   61856: out<=1;
   61857: out<=0;
   61858: out<=0;
   61859: out<=1;
   61860: out<=1;
   61861: out<=1;
   61862: out<=1;
   61863: out<=1;
   61864: out<=1;
   61865: out<=1;
   61866: out<=0;
   61867: out<=0;
   61868: out<=1;
   61869: out<=0;
   61870: out<=1;
   61871: out<=0;
   61872: out<=0;
   61873: out<=0;
   61874: out<=0;
   61875: out<=0;
   61876: out<=1;
   61877: out<=0;
   61878: out<=0;
   61879: out<=1;
   61880: out<=1;
   61881: out<=0;
   61882: out<=1;
   61883: out<=0;
   61884: out<=0;
   61885: out<=0;
   61886: out<=1;
   61887: out<=1;
   61888: out<=0;
   61889: out<=0;
   61890: out<=1;
   61891: out<=1;
   61892: out<=1;
   61893: out<=0;
   61894: out<=1;
   61895: out<=0;
   61896: out<=0;
   61897: out<=1;
   61898: out<=1;
   61899: out<=0;
   61900: out<=1;
   61901: out<=1;
   61902: out<=1;
   61903: out<=1;
   61904: out<=0;
   61905: out<=1;
   61906: out<=0;
   61907: out<=1;
   61908: out<=0;
   61909: out<=0;
   61910: out<=1;
   61911: out<=1;
   61912: out<=1;
   61913: out<=1;
   61914: out<=1;
   61915: out<=1;
   61916: out<=1;
   61917: out<=0;
   61918: out<=0;
   61919: out<=1;
   61920: out<=0;
   61921: out<=1;
   61922: out<=1;
   61923: out<=0;
   61924: out<=0;
   61925: out<=0;
   61926: out<=0;
   61927: out<=0;
   61928: out<=0;
   61929: out<=0;
   61930: out<=1;
   61931: out<=1;
   61932: out<=0;
   61933: out<=1;
   61934: out<=0;
   61935: out<=1;
   61936: out<=0;
   61937: out<=0;
   61938: out<=0;
   61939: out<=0;
   61940: out<=1;
   61941: out<=0;
   61942: out<=0;
   61943: out<=1;
   61944: out<=1;
   61945: out<=0;
   61946: out<=1;
   61947: out<=0;
   61948: out<=0;
   61949: out<=0;
   61950: out<=1;
   61951: out<=1;
   61952: out<=0;
   61953: out<=0;
   61954: out<=0;
   61955: out<=0;
   61956: out<=1;
   61957: out<=0;
   61958: out<=0;
   61959: out<=1;
   61960: out<=1;
   61961: out<=0;
   61962: out<=1;
   61963: out<=0;
   61964: out<=0;
   61965: out<=0;
   61966: out<=1;
   61967: out<=1;
   61968: out<=0;
   61969: out<=1;
   61970: out<=1;
   61971: out<=0;
   61972: out<=0;
   61973: out<=0;
   61974: out<=0;
   61975: out<=0;
   61976: out<=0;
   61977: out<=0;
   61978: out<=1;
   61979: out<=1;
   61980: out<=0;
   61981: out<=1;
   61982: out<=0;
   61983: out<=1;
   61984: out<=0;
   61985: out<=1;
   61986: out<=0;
   61987: out<=1;
   61988: out<=0;
   61989: out<=0;
   61990: out<=1;
   61991: out<=1;
   61992: out<=1;
   61993: out<=1;
   61994: out<=1;
   61995: out<=1;
   61996: out<=1;
   61997: out<=0;
   61998: out<=0;
   61999: out<=1;
   62000: out<=0;
   62001: out<=0;
   62002: out<=1;
   62003: out<=1;
   62004: out<=1;
   62005: out<=0;
   62006: out<=1;
   62007: out<=0;
   62008: out<=0;
   62009: out<=1;
   62010: out<=1;
   62011: out<=0;
   62012: out<=1;
   62013: out<=1;
   62014: out<=1;
   62015: out<=1;
   62016: out<=0;
   62017: out<=0;
   62018: out<=0;
   62019: out<=0;
   62020: out<=1;
   62021: out<=0;
   62022: out<=0;
   62023: out<=1;
   62024: out<=1;
   62025: out<=0;
   62026: out<=1;
   62027: out<=0;
   62028: out<=0;
   62029: out<=0;
   62030: out<=1;
   62031: out<=1;
   62032: out<=1;
   62033: out<=0;
   62034: out<=0;
   62035: out<=1;
   62036: out<=1;
   62037: out<=1;
   62038: out<=1;
   62039: out<=1;
   62040: out<=1;
   62041: out<=1;
   62042: out<=0;
   62043: out<=0;
   62044: out<=1;
   62045: out<=0;
   62046: out<=1;
   62047: out<=0;
   62048: out<=1;
   62049: out<=0;
   62050: out<=1;
   62051: out<=0;
   62052: out<=1;
   62053: out<=1;
   62054: out<=0;
   62055: out<=0;
   62056: out<=0;
   62057: out<=0;
   62058: out<=0;
   62059: out<=0;
   62060: out<=0;
   62061: out<=1;
   62062: out<=1;
   62063: out<=0;
   62064: out<=0;
   62065: out<=0;
   62066: out<=1;
   62067: out<=1;
   62068: out<=1;
   62069: out<=0;
   62070: out<=1;
   62071: out<=0;
   62072: out<=0;
   62073: out<=1;
   62074: out<=1;
   62075: out<=0;
   62076: out<=1;
   62077: out<=1;
   62078: out<=1;
   62079: out<=1;
   62080: out<=1;
   62081: out<=1;
   62082: out<=1;
   62083: out<=1;
   62084: out<=0;
   62085: out<=1;
   62086: out<=1;
   62087: out<=0;
   62088: out<=0;
   62089: out<=1;
   62090: out<=0;
   62091: out<=1;
   62092: out<=1;
   62093: out<=1;
   62094: out<=0;
   62095: out<=0;
   62096: out<=0;
   62097: out<=1;
   62098: out<=1;
   62099: out<=0;
   62100: out<=0;
   62101: out<=0;
   62102: out<=0;
   62103: out<=0;
   62104: out<=0;
   62105: out<=0;
   62106: out<=1;
   62107: out<=1;
   62108: out<=0;
   62109: out<=1;
   62110: out<=0;
   62111: out<=1;
   62112: out<=1;
   62113: out<=0;
   62114: out<=1;
   62115: out<=0;
   62116: out<=1;
   62117: out<=1;
   62118: out<=0;
   62119: out<=0;
   62120: out<=0;
   62121: out<=0;
   62122: out<=0;
   62123: out<=0;
   62124: out<=0;
   62125: out<=1;
   62126: out<=1;
   62127: out<=0;
   62128: out<=0;
   62129: out<=0;
   62130: out<=1;
   62131: out<=1;
   62132: out<=1;
   62133: out<=0;
   62134: out<=1;
   62135: out<=0;
   62136: out<=0;
   62137: out<=1;
   62138: out<=1;
   62139: out<=0;
   62140: out<=1;
   62141: out<=1;
   62142: out<=1;
   62143: out<=1;
   62144: out<=1;
   62145: out<=1;
   62146: out<=1;
   62147: out<=1;
   62148: out<=0;
   62149: out<=1;
   62150: out<=1;
   62151: out<=0;
   62152: out<=0;
   62153: out<=1;
   62154: out<=0;
   62155: out<=1;
   62156: out<=1;
   62157: out<=1;
   62158: out<=0;
   62159: out<=0;
   62160: out<=1;
   62161: out<=0;
   62162: out<=0;
   62163: out<=1;
   62164: out<=1;
   62165: out<=1;
   62166: out<=1;
   62167: out<=1;
   62168: out<=1;
   62169: out<=1;
   62170: out<=0;
   62171: out<=0;
   62172: out<=1;
   62173: out<=0;
   62174: out<=1;
   62175: out<=0;
   62176: out<=0;
   62177: out<=1;
   62178: out<=0;
   62179: out<=1;
   62180: out<=0;
   62181: out<=0;
   62182: out<=1;
   62183: out<=1;
   62184: out<=1;
   62185: out<=1;
   62186: out<=1;
   62187: out<=1;
   62188: out<=1;
   62189: out<=0;
   62190: out<=0;
   62191: out<=1;
   62192: out<=0;
   62193: out<=0;
   62194: out<=1;
   62195: out<=1;
   62196: out<=1;
   62197: out<=0;
   62198: out<=1;
   62199: out<=0;
   62200: out<=0;
   62201: out<=1;
   62202: out<=1;
   62203: out<=0;
   62204: out<=1;
   62205: out<=1;
   62206: out<=1;
   62207: out<=1;
   62208: out<=1;
   62209: out<=0;
   62210: out<=0;
   62211: out<=1;
   62212: out<=1;
   62213: out<=1;
   62214: out<=1;
   62215: out<=1;
   62216: out<=1;
   62217: out<=1;
   62218: out<=0;
   62219: out<=0;
   62220: out<=1;
   62221: out<=0;
   62222: out<=1;
   62223: out<=0;
   62224: out<=0;
   62225: out<=0;
   62226: out<=0;
   62227: out<=0;
   62228: out<=1;
   62229: out<=0;
   62230: out<=0;
   62231: out<=1;
   62232: out<=1;
   62233: out<=0;
   62234: out<=1;
   62235: out<=0;
   62236: out<=0;
   62237: out<=0;
   62238: out<=1;
   62239: out<=1;
   62240: out<=0;
   62241: out<=0;
   62242: out<=1;
   62243: out<=1;
   62244: out<=1;
   62245: out<=0;
   62246: out<=1;
   62247: out<=0;
   62248: out<=0;
   62249: out<=1;
   62250: out<=1;
   62251: out<=0;
   62252: out<=1;
   62253: out<=1;
   62254: out<=1;
   62255: out<=1;
   62256: out<=1;
   62257: out<=0;
   62258: out<=1;
   62259: out<=0;
   62260: out<=1;
   62261: out<=1;
   62262: out<=0;
   62263: out<=0;
   62264: out<=0;
   62265: out<=0;
   62266: out<=0;
   62267: out<=0;
   62268: out<=0;
   62269: out<=1;
   62270: out<=1;
   62271: out<=0;
   62272: out<=0;
   62273: out<=1;
   62274: out<=1;
   62275: out<=0;
   62276: out<=0;
   62277: out<=0;
   62278: out<=0;
   62279: out<=0;
   62280: out<=0;
   62281: out<=0;
   62282: out<=1;
   62283: out<=1;
   62284: out<=0;
   62285: out<=1;
   62286: out<=0;
   62287: out<=1;
   62288: out<=0;
   62289: out<=0;
   62290: out<=0;
   62291: out<=0;
   62292: out<=1;
   62293: out<=0;
   62294: out<=0;
   62295: out<=1;
   62296: out<=1;
   62297: out<=0;
   62298: out<=1;
   62299: out<=0;
   62300: out<=0;
   62301: out<=0;
   62302: out<=1;
   62303: out<=1;
   62304: out<=0;
   62305: out<=0;
   62306: out<=1;
   62307: out<=1;
   62308: out<=1;
   62309: out<=0;
   62310: out<=1;
   62311: out<=0;
   62312: out<=0;
   62313: out<=1;
   62314: out<=1;
   62315: out<=0;
   62316: out<=1;
   62317: out<=1;
   62318: out<=1;
   62319: out<=1;
   62320: out<=0;
   62321: out<=1;
   62322: out<=0;
   62323: out<=1;
   62324: out<=0;
   62325: out<=0;
   62326: out<=1;
   62327: out<=1;
   62328: out<=1;
   62329: out<=1;
   62330: out<=1;
   62331: out<=1;
   62332: out<=1;
   62333: out<=0;
   62334: out<=0;
   62335: out<=1;
   62336: out<=1;
   62337: out<=0;
   62338: out<=0;
   62339: out<=1;
   62340: out<=1;
   62341: out<=1;
   62342: out<=1;
   62343: out<=1;
   62344: out<=1;
   62345: out<=1;
   62346: out<=0;
   62347: out<=0;
   62348: out<=1;
   62349: out<=0;
   62350: out<=1;
   62351: out<=0;
   62352: out<=1;
   62353: out<=1;
   62354: out<=1;
   62355: out<=1;
   62356: out<=0;
   62357: out<=1;
   62358: out<=1;
   62359: out<=0;
   62360: out<=0;
   62361: out<=1;
   62362: out<=0;
   62363: out<=1;
   62364: out<=1;
   62365: out<=1;
   62366: out<=0;
   62367: out<=0;
   62368: out<=0;
   62369: out<=0;
   62370: out<=1;
   62371: out<=1;
   62372: out<=1;
   62373: out<=0;
   62374: out<=1;
   62375: out<=0;
   62376: out<=0;
   62377: out<=1;
   62378: out<=1;
   62379: out<=0;
   62380: out<=1;
   62381: out<=1;
   62382: out<=1;
   62383: out<=1;
   62384: out<=0;
   62385: out<=1;
   62386: out<=0;
   62387: out<=1;
   62388: out<=0;
   62389: out<=0;
   62390: out<=1;
   62391: out<=1;
   62392: out<=1;
   62393: out<=1;
   62394: out<=1;
   62395: out<=1;
   62396: out<=1;
   62397: out<=0;
   62398: out<=0;
   62399: out<=1;
   62400: out<=0;
   62401: out<=1;
   62402: out<=1;
   62403: out<=0;
   62404: out<=0;
   62405: out<=0;
   62406: out<=0;
   62407: out<=0;
   62408: out<=0;
   62409: out<=0;
   62410: out<=1;
   62411: out<=1;
   62412: out<=0;
   62413: out<=1;
   62414: out<=0;
   62415: out<=1;
   62416: out<=1;
   62417: out<=1;
   62418: out<=1;
   62419: out<=1;
   62420: out<=0;
   62421: out<=1;
   62422: out<=1;
   62423: out<=0;
   62424: out<=0;
   62425: out<=1;
   62426: out<=0;
   62427: out<=1;
   62428: out<=1;
   62429: out<=1;
   62430: out<=0;
   62431: out<=0;
   62432: out<=0;
   62433: out<=0;
   62434: out<=1;
   62435: out<=1;
   62436: out<=1;
   62437: out<=0;
   62438: out<=1;
   62439: out<=0;
   62440: out<=0;
   62441: out<=1;
   62442: out<=1;
   62443: out<=0;
   62444: out<=1;
   62445: out<=1;
   62446: out<=1;
   62447: out<=1;
   62448: out<=1;
   62449: out<=0;
   62450: out<=1;
   62451: out<=0;
   62452: out<=1;
   62453: out<=1;
   62454: out<=0;
   62455: out<=0;
   62456: out<=0;
   62457: out<=0;
   62458: out<=0;
   62459: out<=0;
   62460: out<=0;
   62461: out<=1;
   62462: out<=1;
   62463: out<=0;
   62464: out<=0;
   62465: out<=0;
   62466: out<=1;
   62467: out<=1;
   62468: out<=0;
   62469: out<=1;
   62470: out<=0;
   62471: out<=1;
   62472: out<=1;
   62473: out<=0;
   62474: out<=0;
   62475: out<=1;
   62476: out<=1;
   62477: out<=1;
   62478: out<=1;
   62479: out<=1;
   62480: out<=1;
   62481: out<=0;
   62482: out<=1;
   62483: out<=0;
   62484: out<=0;
   62485: out<=0;
   62486: out<=1;
   62487: out<=1;
   62488: out<=1;
   62489: out<=1;
   62490: out<=1;
   62491: out<=1;
   62492: out<=0;
   62493: out<=1;
   62494: out<=1;
   62495: out<=0;
   62496: out<=0;
   62497: out<=1;
   62498: out<=1;
   62499: out<=0;
   62500: out<=1;
   62501: out<=1;
   62502: out<=1;
   62503: out<=1;
   62504: out<=1;
   62505: out<=1;
   62506: out<=0;
   62507: out<=0;
   62508: out<=0;
   62509: out<=1;
   62510: out<=0;
   62511: out<=1;
   62512: out<=1;
   62513: out<=1;
   62514: out<=1;
   62515: out<=1;
   62516: out<=1;
   62517: out<=0;
   62518: out<=0;
   62519: out<=1;
   62520: out<=1;
   62521: out<=0;
   62522: out<=1;
   62523: out<=0;
   62524: out<=1;
   62525: out<=1;
   62526: out<=0;
   62527: out<=0;
   62528: out<=0;
   62529: out<=0;
   62530: out<=1;
   62531: out<=1;
   62532: out<=0;
   62533: out<=1;
   62534: out<=0;
   62535: out<=1;
   62536: out<=1;
   62537: out<=0;
   62538: out<=0;
   62539: out<=1;
   62540: out<=1;
   62541: out<=1;
   62542: out<=1;
   62543: out<=1;
   62544: out<=0;
   62545: out<=1;
   62546: out<=0;
   62547: out<=1;
   62548: out<=1;
   62549: out<=1;
   62550: out<=0;
   62551: out<=0;
   62552: out<=0;
   62553: out<=0;
   62554: out<=0;
   62555: out<=0;
   62556: out<=1;
   62557: out<=0;
   62558: out<=0;
   62559: out<=1;
   62560: out<=1;
   62561: out<=0;
   62562: out<=0;
   62563: out<=1;
   62564: out<=0;
   62565: out<=0;
   62566: out<=0;
   62567: out<=0;
   62568: out<=0;
   62569: out<=0;
   62570: out<=1;
   62571: out<=1;
   62572: out<=1;
   62573: out<=0;
   62574: out<=1;
   62575: out<=0;
   62576: out<=1;
   62577: out<=1;
   62578: out<=1;
   62579: out<=1;
   62580: out<=1;
   62581: out<=0;
   62582: out<=0;
   62583: out<=1;
   62584: out<=1;
   62585: out<=0;
   62586: out<=1;
   62587: out<=0;
   62588: out<=1;
   62589: out<=1;
   62590: out<=0;
   62591: out<=0;
   62592: out<=0;
   62593: out<=0;
   62594: out<=1;
   62595: out<=1;
   62596: out<=0;
   62597: out<=1;
   62598: out<=0;
   62599: out<=1;
   62600: out<=1;
   62601: out<=0;
   62602: out<=0;
   62603: out<=1;
   62604: out<=1;
   62605: out<=1;
   62606: out<=1;
   62607: out<=1;
   62608: out<=0;
   62609: out<=1;
   62610: out<=0;
   62611: out<=1;
   62612: out<=1;
   62613: out<=1;
   62614: out<=0;
   62615: out<=0;
   62616: out<=0;
   62617: out<=0;
   62618: out<=0;
   62619: out<=0;
   62620: out<=1;
   62621: out<=0;
   62622: out<=0;
   62623: out<=1;
   62624: out<=0;
   62625: out<=1;
   62626: out<=1;
   62627: out<=0;
   62628: out<=1;
   62629: out<=1;
   62630: out<=1;
   62631: out<=1;
   62632: out<=1;
   62633: out<=1;
   62634: out<=0;
   62635: out<=0;
   62636: out<=0;
   62637: out<=1;
   62638: out<=0;
   62639: out<=1;
   62640: out<=0;
   62641: out<=0;
   62642: out<=0;
   62643: out<=0;
   62644: out<=0;
   62645: out<=1;
   62646: out<=1;
   62647: out<=0;
   62648: out<=0;
   62649: out<=1;
   62650: out<=0;
   62651: out<=1;
   62652: out<=0;
   62653: out<=0;
   62654: out<=1;
   62655: out<=1;
   62656: out<=0;
   62657: out<=0;
   62658: out<=1;
   62659: out<=1;
   62660: out<=0;
   62661: out<=1;
   62662: out<=0;
   62663: out<=1;
   62664: out<=1;
   62665: out<=0;
   62666: out<=0;
   62667: out<=1;
   62668: out<=1;
   62669: out<=1;
   62670: out<=1;
   62671: out<=1;
   62672: out<=1;
   62673: out<=0;
   62674: out<=1;
   62675: out<=0;
   62676: out<=0;
   62677: out<=0;
   62678: out<=1;
   62679: out<=1;
   62680: out<=1;
   62681: out<=1;
   62682: out<=1;
   62683: out<=1;
   62684: out<=0;
   62685: out<=1;
   62686: out<=1;
   62687: out<=0;
   62688: out<=1;
   62689: out<=0;
   62690: out<=0;
   62691: out<=1;
   62692: out<=0;
   62693: out<=0;
   62694: out<=0;
   62695: out<=0;
   62696: out<=0;
   62697: out<=0;
   62698: out<=1;
   62699: out<=1;
   62700: out<=1;
   62701: out<=0;
   62702: out<=1;
   62703: out<=0;
   62704: out<=0;
   62705: out<=0;
   62706: out<=0;
   62707: out<=0;
   62708: out<=0;
   62709: out<=1;
   62710: out<=1;
   62711: out<=0;
   62712: out<=0;
   62713: out<=1;
   62714: out<=0;
   62715: out<=1;
   62716: out<=0;
   62717: out<=0;
   62718: out<=1;
   62719: out<=1;
   62720: out<=0;
   62721: out<=1;
   62722: out<=0;
   62723: out<=1;
   62724: out<=1;
   62725: out<=1;
   62726: out<=0;
   62727: out<=0;
   62728: out<=0;
   62729: out<=0;
   62730: out<=0;
   62731: out<=0;
   62732: out<=1;
   62733: out<=0;
   62734: out<=0;
   62735: out<=1;
   62736: out<=0;
   62737: out<=0;
   62738: out<=1;
   62739: out<=1;
   62740: out<=0;
   62741: out<=1;
   62742: out<=0;
   62743: out<=1;
   62744: out<=1;
   62745: out<=0;
   62746: out<=0;
   62747: out<=1;
   62748: out<=1;
   62749: out<=1;
   62750: out<=1;
   62751: out<=1;
   62752: out<=1;
   62753: out<=1;
   62754: out<=1;
   62755: out<=1;
   62756: out<=1;
   62757: out<=0;
   62758: out<=0;
   62759: out<=1;
   62760: out<=1;
   62761: out<=0;
   62762: out<=1;
   62763: out<=0;
   62764: out<=1;
   62765: out<=1;
   62766: out<=0;
   62767: out<=0;
   62768: out<=1;
   62769: out<=0;
   62770: out<=0;
   62771: out<=1;
   62772: out<=0;
   62773: out<=0;
   62774: out<=0;
   62775: out<=0;
   62776: out<=0;
   62777: out<=0;
   62778: out<=1;
   62779: out<=1;
   62780: out<=1;
   62781: out<=0;
   62782: out<=1;
   62783: out<=0;
   62784: out<=1;
   62785: out<=0;
   62786: out<=1;
   62787: out<=0;
   62788: out<=0;
   62789: out<=0;
   62790: out<=1;
   62791: out<=1;
   62792: out<=1;
   62793: out<=1;
   62794: out<=1;
   62795: out<=1;
   62796: out<=0;
   62797: out<=1;
   62798: out<=1;
   62799: out<=0;
   62800: out<=0;
   62801: out<=0;
   62802: out<=1;
   62803: out<=1;
   62804: out<=0;
   62805: out<=1;
   62806: out<=0;
   62807: out<=1;
   62808: out<=1;
   62809: out<=0;
   62810: out<=0;
   62811: out<=1;
   62812: out<=1;
   62813: out<=1;
   62814: out<=1;
   62815: out<=1;
   62816: out<=1;
   62817: out<=1;
   62818: out<=1;
   62819: out<=1;
   62820: out<=1;
   62821: out<=0;
   62822: out<=0;
   62823: out<=1;
   62824: out<=1;
   62825: out<=0;
   62826: out<=1;
   62827: out<=0;
   62828: out<=1;
   62829: out<=1;
   62830: out<=0;
   62831: out<=0;
   62832: out<=0;
   62833: out<=1;
   62834: out<=1;
   62835: out<=0;
   62836: out<=1;
   62837: out<=1;
   62838: out<=1;
   62839: out<=1;
   62840: out<=1;
   62841: out<=1;
   62842: out<=0;
   62843: out<=0;
   62844: out<=0;
   62845: out<=1;
   62846: out<=0;
   62847: out<=1;
   62848: out<=1;
   62849: out<=0;
   62850: out<=1;
   62851: out<=0;
   62852: out<=0;
   62853: out<=0;
   62854: out<=1;
   62855: out<=1;
   62856: out<=1;
   62857: out<=1;
   62858: out<=1;
   62859: out<=1;
   62860: out<=0;
   62861: out<=1;
   62862: out<=1;
   62863: out<=0;
   62864: out<=0;
   62865: out<=0;
   62866: out<=1;
   62867: out<=1;
   62868: out<=0;
   62869: out<=1;
   62870: out<=0;
   62871: out<=1;
   62872: out<=1;
   62873: out<=0;
   62874: out<=0;
   62875: out<=1;
   62876: out<=1;
   62877: out<=1;
   62878: out<=1;
   62879: out<=1;
   62880: out<=0;
   62881: out<=0;
   62882: out<=0;
   62883: out<=0;
   62884: out<=0;
   62885: out<=1;
   62886: out<=1;
   62887: out<=0;
   62888: out<=0;
   62889: out<=1;
   62890: out<=0;
   62891: out<=1;
   62892: out<=0;
   62893: out<=0;
   62894: out<=1;
   62895: out<=1;
   62896: out<=1;
   62897: out<=0;
   62898: out<=0;
   62899: out<=1;
   62900: out<=0;
   62901: out<=0;
   62902: out<=0;
   62903: out<=0;
   62904: out<=0;
   62905: out<=0;
   62906: out<=1;
   62907: out<=1;
   62908: out<=1;
   62909: out<=0;
   62910: out<=1;
   62911: out<=0;
   62912: out<=0;
   62913: out<=1;
   62914: out<=0;
   62915: out<=1;
   62916: out<=1;
   62917: out<=1;
   62918: out<=0;
   62919: out<=0;
   62920: out<=0;
   62921: out<=0;
   62922: out<=0;
   62923: out<=0;
   62924: out<=1;
   62925: out<=0;
   62926: out<=0;
   62927: out<=1;
   62928: out<=0;
   62929: out<=0;
   62930: out<=1;
   62931: out<=1;
   62932: out<=0;
   62933: out<=1;
   62934: out<=0;
   62935: out<=1;
   62936: out<=1;
   62937: out<=0;
   62938: out<=0;
   62939: out<=1;
   62940: out<=1;
   62941: out<=1;
   62942: out<=1;
   62943: out<=1;
   62944: out<=0;
   62945: out<=0;
   62946: out<=0;
   62947: out<=0;
   62948: out<=0;
   62949: out<=1;
   62950: out<=1;
   62951: out<=0;
   62952: out<=0;
   62953: out<=1;
   62954: out<=0;
   62955: out<=1;
   62956: out<=0;
   62957: out<=0;
   62958: out<=1;
   62959: out<=1;
   62960: out<=0;
   62961: out<=1;
   62962: out<=1;
   62963: out<=0;
   62964: out<=1;
   62965: out<=1;
   62966: out<=1;
   62967: out<=1;
   62968: out<=1;
   62969: out<=1;
   62970: out<=0;
   62971: out<=0;
   62972: out<=0;
   62973: out<=1;
   62974: out<=0;
   62975: out<=1;
   62976: out<=0;
   62977: out<=1;
   62978: out<=1;
   62979: out<=0;
   62980: out<=1;
   62981: out<=1;
   62982: out<=1;
   62983: out<=1;
   62984: out<=1;
   62985: out<=1;
   62986: out<=0;
   62987: out<=0;
   62988: out<=0;
   62989: out<=1;
   62990: out<=0;
   62991: out<=1;
   62992: out<=0;
   62993: out<=0;
   62994: out<=0;
   62995: out<=0;
   62996: out<=0;
   62997: out<=1;
   62998: out<=1;
   62999: out<=0;
   63000: out<=0;
   63001: out<=1;
   63002: out<=0;
   63003: out<=1;
   63004: out<=0;
   63005: out<=0;
   63006: out<=1;
   63007: out<=1;
   63008: out<=0;
   63009: out<=0;
   63010: out<=1;
   63011: out<=1;
   63012: out<=0;
   63013: out<=1;
   63014: out<=0;
   63015: out<=1;
   63016: out<=1;
   63017: out<=0;
   63018: out<=0;
   63019: out<=1;
   63020: out<=1;
   63021: out<=1;
   63022: out<=1;
   63023: out<=1;
   63024: out<=0;
   63025: out<=1;
   63026: out<=0;
   63027: out<=1;
   63028: out<=1;
   63029: out<=1;
   63030: out<=0;
   63031: out<=0;
   63032: out<=0;
   63033: out<=0;
   63034: out<=0;
   63035: out<=0;
   63036: out<=1;
   63037: out<=0;
   63038: out<=0;
   63039: out<=1;
   63040: out<=1;
   63041: out<=0;
   63042: out<=0;
   63043: out<=1;
   63044: out<=0;
   63045: out<=0;
   63046: out<=0;
   63047: out<=0;
   63048: out<=0;
   63049: out<=0;
   63050: out<=1;
   63051: out<=1;
   63052: out<=1;
   63053: out<=0;
   63054: out<=1;
   63055: out<=0;
   63056: out<=0;
   63057: out<=0;
   63058: out<=0;
   63059: out<=0;
   63060: out<=0;
   63061: out<=1;
   63062: out<=1;
   63063: out<=0;
   63064: out<=0;
   63065: out<=1;
   63066: out<=0;
   63067: out<=1;
   63068: out<=0;
   63069: out<=0;
   63070: out<=1;
   63071: out<=1;
   63072: out<=0;
   63073: out<=0;
   63074: out<=1;
   63075: out<=1;
   63076: out<=0;
   63077: out<=1;
   63078: out<=0;
   63079: out<=1;
   63080: out<=1;
   63081: out<=0;
   63082: out<=0;
   63083: out<=1;
   63084: out<=1;
   63085: out<=1;
   63086: out<=1;
   63087: out<=1;
   63088: out<=1;
   63089: out<=0;
   63090: out<=1;
   63091: out<=0;
   63092: out<=0;
   63093: out<=0;
   63094: out<=1;
   63095: out<=1;
   63096: out<=1;
   63097: out<=1;
   63098: out<=1;
   63099: out<=1;
   63100: out<=0;
   63101: out<=1;
   63102: out<=1;
   63103: out<=0;
   63104: out<=0;
   63105: out<=1;
   63106: out<=1;
   63107: out<=0;
   63108: out<=1;
   63109: out<=1;
   63110: out<=1;
   63111: out<=1;
   63112: out<=1;
   63113: out<=1;
   63114: out<=0;
   63115: out<=0;
   63116: out<=0;
   63117: out<=1;
   63118: out<=0;
   63119: out<=1;
   63120: out<=1;
   63121: out<=1;
   63122: out<=1;
   63123: out<=1;
   63124: out<=1;
   63125: out<=0;
   63126: out<=0;
   63127: out<=1;
   63128: out<=1;
   63129: out<=0;
   63130: out<=1;
   63131: out<=0;
   63132: out<=1;
   63133: out<=1;
   63134: out<=0;
   63135: out<=0;
   63136: out<=0;
   63137: out<=0;
   63138: out<=1;
   63139: out<=1;
   63140: out<=0;
   63141: out<=1;
   63142: out<=0;
   63143: out<=1;
   63144: out<=1;
   63145: out<=0;
   63146: out<=0;
   63147: out<=1;
   63148: out<=1;
   63149: out<=1;
   63150: out<=1;
   63151: out<=1;
   63152: out<=1;
   63153: out<=0;
   63154: out<=1;
   63155: out<=0;
   63156: out<=0;
   63157: out<=0;
   63158: out<=1;
   63159: out<=1;
   63160: out<=1;
   63161: out<=1;
   63162: out<=1;
   63163: out<=1;
   63164: out<=0;
   63165: out<=1;
   63166: out<=1;
   63167: out<=0;
   63168: out<=1;
   63169: out<=0;
   63170: out<=0;
   63171: out<=1;
   63172: out<=0;
   63173: out<=0;
   63174: out<=0;
   63175: out<=0;
   63176: out<=0;
   63177: out<=0;
   63178: out<=1;
   63179: out<=1;
   63180: out<=1;
   63181: out<=0;
   63182: out<=1;
   63183: out<=0;
   63184: out<=1;
   63185: out<=1;
   63186: out<=1;
   63187: out<=1;
   63188: out<=1;
   63189: out<=0;
   63190: out<=0;
   63191: out<=1;
   63192: out<=1;
   63193: out<=0;
   63194: out<=1;
   63195: out<=0;
   63196: out<=1;
   63197: out<=1;
   63198: out<=0;
   63199: out<=0;
   63200: out<=0;
   63201: out<=0;
   63202: out<=1;
   63203: out<=1;
   63204: out<=0;
   63205: out<=1;
   63206: out<=0;
   63207: out<=1;
   63208: out<=1;
   63209: out<=0;
   63210: out<=0;
   63211: out<=1;
   63212: out<=1;
   63213: out<=1;
   63214: out<=1;
   63215: out<=1;
   63216: out<=0;
   63217: out<=1;
   63218: out<=0;
   63219: out<=1;
   63220: out<=1;
   63221: out<=1;
   63222: out<=0;
   63223: out<=0;
   63224: out<=0;
   63225: out<=0;
   63226: out<=0;
   63227: out<=0;
   63228: out<=1;
   63229: out<=0;
   63230: out<=0;
   63231: out<=1;
   63232: out<=0;
   63233: out<=0;
   63234: out<=0;
   63235: out<=0;
   63236: out<=0;
   63237: out<=1;
   63238: out<=1;
   63239: out<=0;
   63240: out<=0;
   63241: out<=1;
   63242: out<=0;
   63243: out<=1;
   63244: out<=0;
   63245: out<=0;
   63246: out<=1;
   63247: out<=1;
   63248: out<=1;
   63249: out<=0;
   63250: out<=0;
   63251: out<=1;
   63252: out<=0;
   63253: out<=0;
   63254: out<=0;
   63255: out<=0;
   63256: out<=0;
   63257: out<=0;
   63258: out<=1;
   63259: out<=1;
   63260: out<=1;
   63261: out<=0;
   63262: out<=1;
   63263: out<=0;
   63264: out<=1;
   63265: out<=0;
   63266: out<=1;
   63267: out<=0;
   63268: out<=0;
   63269: out<=0;
   63270: out<=1;
   63271: out<=1;
   63272: out<=1;
   63273: out<=1;
   63274: out<=1;
   63275: out<=1;
   63276: out<=0;
   63277: out<=1;
   63278: out<=1;
   63279: out<=0;
   63280: out<=0;
   63281: out<=0;
   63282: out<=1;
   63283: out<=1;
   63284: out<=0;
   63285: out<=1;
   63286: out<=0;
   63287: out<=1;
   63288: out<=1;
   63289: out<=0;
   63290: out<=0;
   63291: out<=1;
   63292: out<=1;
   63293: out<=1;
   63294: out<=1;
   63295: out<=1;
   63296: out<=0;
   63297: out<=0;
   63298: out<=0;
   63299: out<=0;
   63300: out<=0;
   63301: out<=1;
   63302: out<=1;
   63303: out<=0;
   63304: out<=0;
   63305: out<=1;
   63306: out<=0;
   63307: out<=1;
   63308: out<=0;
   63309: out<=0;
   63310: out<=1;
   63311: out<=1;
   63312: out<=0;
   63313: out<=1;
   63314: out<=1;
   63315: out<=0;
   63316: out<=1;
   63317: out<=1;
   63318: out<=1;
   63319: out<=1;
   63320: out<=1;
   63321: out<=1;
   63322: out<=0;
   63323: out<=0;
   63324: out<=0;
   63325: out<=1;
   63326: out<=0;
   63327: out<=1;
   63328: out<=0;
   63329: out<=1;
   63330: out<=0;
   63331: out<=1;
   63332: out<=1;
   63333: out<=1;
   63334: out<=0;
   63335: out<=0;
   63336: out<=0;
   63337: out<=0;
   63338: out<=0;
   63339: out<=0;
   63340: out<=1;
   63341: out<=0;
   63342: out<=0;
   63343: out<=1;
   63344: out<=0;
   63345: out<=0;
   63346: out<=1;
   63347: out<=1;
   63348: out<=0;
   63349: out<=1;
   63350: out<=0;
   63351: out<=1;
   63352: out<=1;
   63353: out<=0;
   63354: out<=0;
   63355: out<=1;
   63356: out<=1;
   63357: out<=1;
   63358: out<=1;
   63359: out<=1;
   63360: out<=1;
   63361: out<=1;
   63362: out<=1;
   63363: out<=1;
   63364: out<=1;
   63365: out<=0;
   63366: out<=0;
   63367: out<=1;
   63368: out<=1;
   63369: out<=0;
   63370: out<=1;
   63371: out<=0;
   63372: out<=1;
   63373: out<=1;
   63374: out<=0;
   63375: out<=0;
   63376: out<=1;
   63377: out<=0;
   63378: out<=0;
   63379: out<=1;
   63380: out<=0;
   63381: out<=0;
   63382: out<=0;
   63383: out<=0;
   63384: out<=0;
   63385: out<=0;
   63386: out<=1;
   63387: out<=1;
   63388: out<=1;
   63389: out<=0;
   63390: out<=1;
   63391: out<=0;
   63392: out<=0;
   63393: out<=1;
   63394: out<=0;
   63395: out<=1;
   63396: out<=1;
   63397: out<=1;
   63398: out<=0;
   63399: out<=0;
   63400: out<=0;
   63401: out<=0;
   63402: out<=0;
   63403: out<=0;
   63404: out<=1;
   63405: out<=0;
   63406: out<=0;
   63407: out<=1;
   63408: out<=0;
   63409: out<=0;
   63410: out<=1;
   63411: out<=1;
   63412: out<=0;
   63413: out<=1;
   63414: out<=0;
   63415: out<=1;
   63416: out<=1;
   63417: out<=0;
   63418: out<=0;
   63419: out<=1;
   63420: out<=1;
   63421: out<=1;
   63422: out<=1;
   63423: out<=1;
   63424: out<=1;
   63425: out<=1;
   63426: out<=1;
   63427: out<=1;
   63428: out<=1;
   63429: out<=0;
   63430: out<=0;
   63431: out<=1;
   63432: out<=1;
   63433: out<=0;
   63434: out<=1;
   63435: out<=0;
   63436: out<=1;
   63437: out<=1;
   63438: out<=0;
   63439: out<=0;
   63440: out<=0;
   63441: out<=1;
   63442: out<=1;
   63443: out<=0;
   63444: out<=1;
   63445: out<=1;
   63446: out<=1;
   63447: out<=1;
   63448: out<=1;
   63449: out<=1;
   63450: out<=0;
   63451: out<=0;
   63452: out<=0;
   63453: out<=1;
   63454: out<=0;
   63455: out<=1;
   63456: out<=1;
   63457: out<=0;
   63458: out<=1;
   63459: out<=0;
   63460: out<=0;
   63461: out<=0;
   63462: out<=1;
   63463: out<=1;
   63464: out<=1;
   63465: out<=1;
   63466: out<=1;
   63467: out<=1;
   63468: out<=0;
   63469: out<=1;
   63470: out<=1;
   63471: out<=0;
   63472: out<=0;
   63473: out<=0;
   63474: out<=1;
   63475: out<=1;
   63476: out<=0;
   63477: out<=1;
   63478: out<=0;
   63479: out<=1;
   63480: out<=1;
   63481: out<=0;
   63482: out<=0;
   63483: out<=1;
   63484: out<=1;
   63485: out<=1;
   63486: out<=1;
   63487: out<=1;
   63488: out<=0;
   63489: out<=0;
   63490: out<=0;
   63491: out<=0;
   63492: out<=0;
   63493: out<=1;
   63494: out<=1;
   63495: out<=0;
   63496: out<=1;
   63497: out<=0;
   63498: out<=1;
   63499: out<=0;
   63500: out<=1;
   63501: out<=1;
   63502: out<=0;
   63503: out<=0;
   63504: out<=1;
   63505: out<=0;
   63506: out<=0;
   63507: out<=1;
   63508: out<=0;
   63509: out<=0;
   63510: out<=0;
   63511: out<=0;
   63512: out<=1;
   63513: out<=1;
   63514: out<=0;
   63515: out<=0;
   63516: out<=0;
   63517: out<=1;
   63518: out<=0;
   63519: out<=1;
   63520: out<=0;
   63521: out<=1;
   63522: out<=0;
   63523: out<=1;
   63524: out<=1;
   63525: out<=1;
   63526: out<=0;
   63527: out<=0;
   63528: out<=1;
   63529: out<=1;
   63530: out<=1;
   63531: out<=1;
   63532: out<=0;
   63533: out<=1;
   63534: out<=1;
   63535: out<=0;
   63536: out<=1;
   63537: out<=1;
   63538: out<=0;
   63539: out<=0;
   63540: out<=1;
   63541: out<=0;
   63542: out<=1;
   63543: out<=0;
   63544: out<=1;
   63545: out<=0;
   63546: out<=0;
   63547: out<=1;
   63548: out<=1;
   63549: out<=1;
   63550: out<=1;
   63551: out<=1;
   63552: out<=0;
   63553: out<=0;
   63554: out<=0;
   63555: out<=0;
   63556: out<=0;
   63557: out<=1;
   63558: out<=1;
   63559: out<=0;
   63560: out<=1;
   63561: out<=0;
   63562: out<=1;
   63563: out<=0;
   63564: out<=1;
   63565: out<=1;
   63566: out<=0;
   63567: out<=0;
   63568: out<=0;
   63569: out<=1;
   63570: out<=1;
   63571: out<=0;
   63572: out<=1;
   63573: out<=1;
   63574: out<=1;
   63575: out<=1;
   63576: out<=0;
   63577: out<=0;
   63578: out<=1;
   63579: out<=1;
   63580: out<=1;
   63581: out<=0;
   63582: out<=1;
   63583: out<=0;
   63584: out<=1;
   63585: out<=0;
   63586: out<=1;
   63587: out<=0;
   63588: out<=0;
   63589: out<=0;
   63590: out<=1;
   63591: out<=1;
   63592: out<=0;
   63593: out<=0;
   63594: out<=0;
   63595: out<=0;
   63596: out<=1;
   63597: out<=0;
   63598: out<=0;
   63599: out<=1;
   63600: out<=1;
   63601: out<=1;
   63602: out<=0;
   63603: out<=0;
   63604: out<=1;
   63605: out<=0;
   63606: out<=1;
   63607: out<=0;
   63608: out<=1;
   63609: out<=0;
   63610: out<=0;
   63611: out<=1;
   63612: out<=1;
   63613: out<=1;
   63614: out<=1;
   63615: out<=1;
   63616: out<=1;
   63617: out<=1;
   63618: out<=1;
   63619: out<=1;
   63620: out<=1;
   63621: out<=0;
   63622: out<=0;
   63623: out<=1;
   63624: out<=0;
   63625: out<=1;
   63626: out<=0;
   63627: out<=1;
   63628: out<=0;
   63629: out<=0;
   63630: out<=1;
   63631: out<=1;
   63632: out<=1;
   63633: out<=0;
   63634: out<=0;
   63635: out<=1;
   63636: out<=0;
   63637: out<=0;
   63638: out<=0;
   63639: out<=0;
   63640: out<=1;
   63641: out<=1;
   63642: out<=0;
   63643: out<=0;
   63644: out<=0;
   63645: out<=1;
   63646: out<=0;
   63647: out<=1;
   63648: out<=1;
   63649: out<=0;
   63650: out<=1;
   63651: out<=0;
   63652: out<=0;
   63653: out<=0;
   63654: out<=1;
   63655: out<=1;
   63656: out<=0;
   63657: out<=0;
   63658: out<=0;
   63659: out<=0;
   63660: out<=1;
   63661: out<=0;
   63662: out<=0;
   63663: out<=1;
   63664: out<=1;
   63665: out<=1;
   63666: out<=0;
   63667: out<=0;
   63668: out<=1;
   63669: out<=0;
   63670: out<=1;
   63671: out<=0;
   63672: out<=1;
   63673: out<=0;
   63674: out<=0;
   63675: out<=1;
   63676: out<=1;
   63677: out<=1;
   63678: out<=1;
   63679: out<=1;
   63680: out<=1;
   63681: out<=1;
   63682: out<=1;
   63683: out<=1;
   63684: out<=1;
   63685: out<=0;
   63686: out<=0;
   63687: out<=1;
   63688: out<=0;
   63689: out<=1;
   63690: out<=0;
   63691: out<=1;
   63692: out<=0;
   63693: out<=0;
   63694: out<=1;
   63695: out<=1;
   63696: out<=0;
   63697: out<=1;
   63698: out<=1;
   63699: out<=0;
   63700: out<=1;
   63701: out<=1;
   63702: out<=1;
   63703: out<=1;
   63704: out<=0;
   63705: out<=0;
   63706: out<=1;
   63707: out<=1;
   63708: out<=1;
   63709: out<=0;
   63710: out<=1;
   63711: out<=0;
   63712: out<=0;
   63713: out<=1;
   63714: out<=0;
   63715: out<=1;
   63716: out<=1;
   63717: out<=1;
   63718: out<=0;
   63719: out<=0;
   63720: out<=1;
   63721: out<=1;
   63722: out<=1;
   63723: out<=1;
   63724: out<=0;
   63725: out<=1;
   63726: out<=1;
   63727: out<=0;
   63728: out<=1;
   63729: out<=1;
   63730: out<=0;
   63731: out<=0;
   63732: out<=1;
   63733: out<=0;
   63734: out<=1;
   63735: out<=0;
   63736: out<=1;
   63737: out<=0;
   63738: out<=0;
   63739: out<=1;
   63740: out<=1;
   63741: out<=1;
   63742: out<=1;
   63743: out<=1;
   63744: out<=0;
   63745: out<=1;
   63746: out<=1;
   63747: out<=0;
   63748: out<=1;
   63749: out<=1;
   63750: out<=1;
   63751: out<=1;
   63752: out<=0;
   63753: out<=0;
   63754: out<=1;
   63755: out<=1;
   63756: out<=1;
   63757: out<=0;
   63758: out<=1;
   63759: out<=0;
   63760: out<=0;
   63761: out<=0;
   63762: out<=0;
   63763: out<=0;
   63764: out<=0;
   63765: out<=1;
   63766: out<=1;
   63767: out<=0;
   63768: out<=1;
   63769: out<=0;
   63770: out<=1;
   63771: out<=0;
   63772: out<=1;
   63773: out<=1;
   63774: out<=0;
   63775: out<=0;
   63776: out<=1;
   63777: out<=1;
   63778: out<=0;
   63779: out<=0;
   63780: out<=1;
   63781: out<=0;
   63782: out<=1;
   63783: out<=0;
   63784: out<=1;
   63785: out<=0;
   63786: out<=0;
   63787: out<=1;
   63788: out<=1;
   63789: out<=1;
   63790: out<=1;
   63791: out<=1;
   63792: out<=1;
   63793: out<=0;
   63794: out<=1;
   63795: out<=0;
   63796: out<=0;
   63797: out<=0;
   63798: out<=1;
   63799: out<=1;
   63800: out<=0;
   63801: out<=0;
   63802: out<=0;
   63803: out<=0;
   63804: out<=1;
   63805: out<=0;
   63806: out<=0;
   63807: out<=1;
   63808: out<=1;
   63809: out<=0;
   63810: out<=0;
   63811: out<=1;
   63812: out<=0;
   63813: out<=0;
   63814: out<=0;
   63815: out<=0;
   63816: out<=1;
   63817: out<=1;
   63818: out<=0;
   63819: out<=0;
   63820: out<=0;
   63821: out<=1;
   63822: out<=0;
   63823: out<=1;
   63824: out<=0;
   63825: out<=0;
   63826: out<=0;
   63827: out<=0;
   63828: out<=0;
   63829: out<=1;
   63830: out<=1;
   63831: out<=0;
   63832: out<=1;
   63833: out<=0;
   63834: out<=1;
   63835: out<=0;
   63836: out<=1;
   63837: out<=1;
   63838: out<=0;
   63839: out<=0;
   63840: out<=1;
   63841: out<=1;
   63842: out<=0;
   63843: out<=0;
   63844: out<=1;
   63845: out<=0;
   63846: out<=1;
   63847: out<=0;
   63848: out<=1;
   63849: out<=0;
   63850: out<=0;
   63851: out<=1;
   63852: out<=1;
   63853: out<=1;
   63854: out<=1;
   63855: out<=1;
   63856: out<=0;
   63857: out<=1;
   63858: out<=0;
   63859: out<=1;
   63860: out<=1;
   63861: out<=1;
   63862: out<=0;
   63863: out<=0;
   63864: out<=1;
   63865: out<=1;
   63866: out<=1;
   63867: out<=1;
   63868: out<=0;
   63869: out<=1;
   63870: out<=1;
   63871: out<=0;
   63872: out<=0;
   63873: out<=1;
   63874: out<=1;
   63875: out<=0;
   63876: out<=1;
   63877: out<=1;
   63878: out<=1;
   63879: out<=1;
   63880: out<=0;
   63881: out<=0;
   63882: out<=1;
   63883: out<=1;
   63884: out<=1;
   63885: out<=0;
   63886: out<=1;
   63887: out<=0;
   63888: out<=1;
   63889: out<=1;
   63890: out<=1;
   63891: out<=1;
   63892: out<=1;
   63893: out<=0;
   63894: out<=0;
   63895: out<=1;
   63896: out<=0;
   63897: out<=1;
   63898: out<=0;
   63899: out<=1;
   63900: out<=0;
   63901: out<=0;
   63902: out<=1;
   63903: out<=1;
   63904: out<=1;
   63905: out<=1;
   63906: out<=0;
   63907: out<=0;
   63908: out<=1;
   63909: out<=0;
   63910: out<=1;
   63911: out<=0;
   63912: out<=1;
   63913: out<=0;
   63914: out<=0;
   63915: out<=1;
   63916: out<=1;
   63917: out<=1;
   63918: out<=1;
   63919: out<=1;
   63920: out<=0;
   63921: out<=1;
   63922: out<=0;
   63923: out<=1;
   63924: out<=1;
   63925: out<=1;
   63926: out<=0;
   63927: out<=0;
   63928: out<=1;
   63929: out<=1;
   63930: out<=1;
   63931: out<=1;
   63932: out<=0;
   63933: out<=1;
   63934: out<=1;
   63935: out<=0;
   63936: out<=1;
   63937: out<=0;
   63938: out<=0;
   63939: out<=1;
   63940: out<=0;
   63941: out<=0;
   63942: out<=0;
   63943: out<=0;
   63944: out<=1;
   63945: out<=1;
   63946: out<=0;
   63947: out<=0;
   63948: out<=0;
   63949: out<=1;
   63950: out<=0;
   63951: out<=1;
   63952: out<=1;
   63953: out<=1;
   63954: out<=1;
   63955: out<=1;
   63956: out<=1;
   63957: out<=0;
   63958: out<=0;
   63959: out<=1;
   63960: out<=0;
   63961: out<=1;
   63962: out<=0;
   63963: out<=1;
   63964: out<=0;
   63965: out<=0;
   63966: out<=1;
   63967: out<=1;
   63968: out<=1;
   63969: out<=1;
   63970: out<=0;
   63971: out<=0;
   63972: out<=1;
   63973: out<=0;
   63974: out<=1;
   63975: out<=0;
   63976: out<=1;
   63977: out<=0;
   63978: out<=0;
   63979: out<=1;
   63980: out<=1;
   63981: out<=1;
   63982: out<=1;
   63983: out<=1;
   63984: out<=1;
   63985: out<=0;
   63986: out<=1;
   63987: out<=0;
   63988: out<=0;
   63989: out<=0;
   63990: out<=1;
   63991: out<=1;
   63992: out<=0;
   63993: out<=0;
   63994: out<=0;
   63995: out<=0;
   63996: out<=1;
   63997: out<=0;
   63998: out<=0;
   63999: out<=1;
   64000: out<=1;
   64001: out<=0;
   64002: out<=1;
   64003: out<=0;
   64004: out<=0;
   64005: out<=0;
   64006: out<=1;
   64007: out<=1;
   64008: out<=0;
   64009: out<=0;
   64010: out<=0;
   64011: out<=0;
   64012: out<=1;
   64013: out<=0;
   64014: out<=0;
   64015: out<=1;
   64016: out<=1;
   64017: out<=1;
   64018: out<=0;
   64019: out<=0;
   64020: out<=1;
   64021: out<=0;
   64022: out<=1;
   64023: out<=0;
   64024: out<=1;
   64025: out<=0;
   64026: out<=0;
   64027: out<=1;
   64028: out<=1;
   64029: out<=1;
   64030: out<=1;
   64031: out<=1;
   64032: out<=1;
   64033: out<=1;
   64034: out<=1;
   64035: out<=1;
   64036: out<=1;
   64037: out<=0;
   64038: out<=0;
   64039: out<=1;
   64040: out<=0;
   64041: out<=1;
   64042: out<=0;
   64043: out<=1;
   64044: out<=0;
   64045: out<=0;
   64046: out<=1;
   64047: out<=1;
   64048: out<=1;
   64049: out<=0;
   64050: out<=0;
   64051: out<=1;
   64052: out<=0;
   64053: out<=0;
   64054: out<=0;
   64055: out<=0;
   64056: out<=1;
   64057: out<=1;
   64058: out<=0;
   64059: out<=0;
   64060: out<=0;
   64061: out<=1;
   64062: out<=0;
   64063: out<=1;
   64064: out<=0;
   64065: out<=1;
   64066: out<=0;
   64067: out<=1;
   64068: out<=1;
   64069: out<=1;
   64070: out<=0;
   64071: out<=0;
   64072: out<=1;
   64073: out<=1;
   64074: out<=1;
   64075: out<=1;
   64076: out<=0;
   64077: out<=1;
   64078: out<=1;
   64079: out<=0;
   64080: out<=1;
   64081: out<=1;
   64082: out<=0;
   64083: out<=0;
   64084: out<=1;
   64085: out<=0;
   64086: out<=1;
   64087: out<=0;
   64088: out<=1;
   64089: out<=0;
   64090: out<=0;
   64091: out<=1;
   64092: out<=1;
   64093: out<=1;
   64094: out<=1;
   64095: out<=1;
   64096: out<=1;
   64097: out<=1;
   64098: out<=1;
   64099: out<=1;
   64100: out<=1;
   64101: out<=0;
   64102: out<=0;
   64103: out<=1;
   64104: out<=0;
   64105: out<=1;
   64106: out<=0;
   64107: out<=1;
   64108: out<=0;
   64109: out<=0;
   64110: out<=1;
   64111: out<=1;
   64112: out<=0;
   64113: out<=1;
   64114: out<=1;
   64115: out<=0;
   64116: out<=1;
   64117: out<=1;
   64118: out<=1;
   64119: out<=1;
   64120: out<=0;
   64121: out<=0;
   64122: out<=1;
   64123: out<=1;
   64124: out<=1;
   64125: out<=0;
   64126: out<=1;
   64127: out<=0;
   64128: out<=0;
   64129: out<=1;
   64130: out<=0;
   64131: out<=1;
   64132: out<=1;
   64133: out<=1;
   64134: out<=0;
   64135: out<=0;
   64136: out<=1;
   64137: out<=1;
   64138: out<=1;
   64139: out<=1;
   64140: out<=0;
   64141: out<=1;
   64142: out<=1;
   64143: out<=0;
   64144: out<=1;
   64145: out<=1;
   64146: out<=0;
   64147: out<=0;
   64148: out<=1;
   64149: out<=0;
   64150: out<=1;
   64151: out<=0;
   64152: out<=1;
   64153: out<=0;
   64154: out<=0;
   64155: out<=1;
   64156: out<=1;
   64157: out<=1;
   64158: out<=1;
   64159: out<=1;
   64160: out<=0;
   64161: out<=0;
   64162: out<=0;
   64163: out<=0;
   64164: out<=0;
   64165: out<=1;
   64166: out<=1;
   64167: out<=0;
   64168: out<=1;
   64169: out<=0;
   64170: out<=1;
   64171: out<=0;
   64172: out<=1;
   64173: out<=1;
   64174: out<=0;
   64175: out<=0;
   64176: out<=1;
   64177: out<=0;
   64178: out<=0;
   64179: out<=1;
   64180: out<=0;
   64181: out<=0;
   64182: out<=0;
   64183: out<=0;
   64184: out<=1;
   64185: out<=1;
   64186: out<=0;
   64187: out<=0;
   64188: out<=0;
   64189: out<=1;
   64190: out<=0;
   64191: out<=1;
   64192: out<=1;
   64193: out<=0;
   64194: out<=1;
   64195: out<=0;
   64196: out<=0;
   64197: out<=0;
   64198: out<=1;
   64199: out<=1;
   64200: out<=0;
   64201: out<=0;
   64202: out<=0;
   64203: out<=0;
   64204: out<=1;
   64205: out<=0;
   64206: out<=0;
   64207: out<=1;
   64208: out<=1;
   64209: out<=1;
   64210: out<=0;
   64211: out<=0;
   64212: out<=1;
   64213: out<=0;
   64214: out<=1;
   64215: out<=0;
   64216: out<=1;
   64217: out<=0;
   64218: out<=0;
   64219: out<=1;
   64220: out<=1;
   64221: out<=1;
   64222: out<=1;
   64223: out<=1;
   64224: out<=0;
   64225: out<=0;
   64226: out<=0;
   64227: out<=0;
   64228: out<=0;
   64229: out<=1;
   64230: out<=1;
   64231: out<=0;
   64232: out<=1;
   64233: out<=0;
   64234: out<=1;
   64235: out<=0;
   64236: out<=1;
   64237: out<=1;
   64238: out<=0;
   64239: out<=0;
   64240: out<=0;
   64241: out<=1;
   64242: out<=1;
   64243: out<=0;
   64244: out<=1;
   64245: out<=1;
   64246: out<=1;
   64247: out<=1;
   64248: out<=0;
   64249: out<=0;
   64250: out<=1;
   64251: out<=1;
   64252: out<=1;
   64253: out<=0;
   64254: out<=1;
   64255: out<=0;
   64256: out<=1;
   64257: out<=1;
   64258: out<=0;
   64259: out<=0;
   64260: out<=1;
   64261: out<=0;
   64262: out<=1;
   64263: out<=0;
   64264: out<=1;
   64265: out<=0;
   64266: out<=0;
   64267: out<=1;
   64268: out<=1;
   64269: out<=1;
   64270: out<=1;
   64271: out<=1;
   64272: out<=0;
   64273: out<=1;
   64274: out<=0;
   64275: out<=1;
   64276: out<=1;
   64277: out<=1;
   64278: out<=0;
   64279: out<=0;
   64280: out<=1;
   64281: out<=1;
   64282: out<=1;
   64283: out<=1;
   64284: out<=0;
   64285: out<=1;
   64286: out<=1;
   64287: out<=0;
   64288: out<=0;
   64289: out<=1;
   64290: out<=1;
   64291: out<=0;
   64292: out<=1;
   64293: out<=1;
   64294: out<=1;
   64295: out<=1;
   64296: out<=0;
   64297: out<=0;
   64298: out<=1;
   64299: out<=1;
   64300: out<=1;
   64301: out<=0;
   64302: out<=1;
   64303: out<=0;
   64304: out<=1;
   64305: out<=1;
   64306: out<=1;
   64307: out<=1;
   64308: out<=1;
   64309: out<=0;
   64310: out<=0;
   64311: out<=1;
   64312: out<=0;
   64313: out<=1;
   64314: out<=0;
   64315: out<=1;
   64316: out<=0;
   64317: out<=0;
   64318: out<=1;
   64319: out<=1;
   64320: out<=1;
   64321: out<=1;
   64322: out<=0;
   64323: out<=0;
   64324: out<=1;
   64325: out<=0;
   64326: out<=1;
   64327: out<=0;
   64328: out<=1;
   64329: out<=0;
   64330: out<=0;
   64331: out<=1;
   64332: out<=1;
   64333: out<=1;
   64334: out<=1;
   64335: out<=1;
   64336: out<=1;
   64337: out<=0;
   64338: out<=1;
   64339: out<=0;
   64340: out<=0;
   64341: out<=0;
   64342: out<=1;
   64343: out<=1;
   64344: out<=0;
   64345: out<=0;
   64346: out<=0;
   64347: out<=0;
   64348: out<=1;
   64349: out<=0;
   64350: out<=0;
   64351: out<=1;
   64352: out<=1;
   64353: out<=0;
   64354: out<=0;
   64355: out<=1;
   64356: out<=0;
   64357: out<=0;
   64358: out<=0;
   64359: out<=0;
   64360: out<=1;
   64361: out<=1;
   64362: out<=0;
   64363: out<=0;
   64364: out<=0;
   64365: out<=1;
   64366: out<=0;
   64367: out<=1;
   64368: out<=1;
   64369: out<=1;
   64370: out<=1;
   64371: out<=1;
   64372: out<=1;
   64373: out<=0;
   64374: out<=0;
   64375: out<=1;
   64376: out<=0;
   64377: out<=1;
   64378: out<=0;
   64379: out<=1;
   64380: out<=0;
   64381: out<=0;
   64382: out<=1;
   64383: out<=1;
   64384: out<=1;
   64385: out<=1;
   64386: out<=0;
   64387: out<=0;
   64388: out<=1;
   64389: out<=0;
   64390: out<=1;
   64391: out<=0;
   64392: out<=1;
   64393: out<=0;
   64394: out<=0;
   64395: out<=1;
   64396: out<=1;
   64397: out<=1;
   64398: out<=1;
   64399: out<=1;
   64400: out<=1;
   64401: out<=0;
   64402: out<=1;
   64403: out<=0;
   64404: out<=0;
   64405: out<=0;
   64406: out<=1;
   64407: out<=1;
   64408: out<=0;
   64409: out<=0;
   64410: out<=0;
   64411: out<=0;
   64412: out<=1;
   64413: out<=0;
   64414: out<=0;
   64415: out<=1;
   64416: out<=0;
   64417: out<=1;
   64418: out<=1;
   64419: out<=0;
   64420: out<=1;
   64421: out<=1;
   64422: out<=1;
   64423: out<=1;
   64424: out<=0;
   64425: out<=0;
   64426: out<=1;
   64427: out<=1;
   64428: out<=1;
   64429: out<=0;
   64430: out<=1;
   64431: out<=0;
   64432: out<=0;
   64433: out<=0;
   64434: out<=0;
   64435: out<=0;
   64436: out<=0;
   64437: out<=1;
   64438: out<=1;
   64439: out<=0;
   64440: out<=1;
   64441: out<=0;
   64442: out<=1;
   64443: out<=0;
   64444: out<=1;
   64445: out<=1;
   64446: out<=0;
   64447: out<=0;
   64448: out<=1;
   64449: out<=1;
   64450: out<=0;
   64451: out<=0;
   64452: out<=1;
   64453: out<=0;
   64454: out<=1;
   64455: out<=0;
   64456: out<=1;
   64457: out<=0;
   64458: out<=0;
   64459: out<=1;
   64460: out<=1;
   64461: out<=1;
   64462: out<=1;
   64463: out<=1;
   64464: out<=0;
   64465: out<=1;
   64466: out<=0;
   64467: out<=1;
   64468: out<=1;
   64469: out<=1;
   64470: out<=0;
   64471: out<=0;
   64472: out<=1;
   64473: out<=1;
   64474: out<=1;
   64475: out<=1;
   64476: out<=0;
   64477: out<=1;
   64478: out<=1;
   64479: out<=0;
   64480: out<=1;
   64481: out<=0;
   64482: out<=0;
   64483: out<=1;
   64484: out<=0;
   64485: out<=0;
   64486: out<=0;
   64487: out<=0;
   64488: out<=1;
   64489: out<=1;
   64490: out<=0;
   64491: out<=0;
   64492: out<=0;
   64493: out<=1;
   64494: out<=0;
   64495: out<=1;
   64496: out<=0;
   64497: out<=0;
   64498: out<=0;
   64499: out<=0;
   64500: out<=0;
   64501: out<=1;
   64502: out<=1;
   64503: out<=0;
   64504: out<=1;
   64505: out<=0;
   64506: out<=1;
   64507: out<=0;
   64508: out<=1;
   64509: out<=1;
   64510: out<=0;
   64511: out<=0;
   64512: out<=1;
   64513: out<=0;
   64514: out<=0;
   64515: out<=1;
   64516: out<=1;
   64517: out<=1;
   64518: out<=1;
   64519: out<=1;
   64520: out<=0;
   64521: out<=0;
   64522: out<=1;
   64523: out<=1;
   64524: out<=0;
   64525: out<=1;
   64526: out<=0;
   64527: out<=1;
   64528: out<=0;
   64529: out<=0;
   64530: out<=0;
   64531: out<=0;
   64532: out<=1;
   64533: out<=0;
   64534: out<=0;
   64535: out<=1;
   64536: out<=0;
   64537: out<=1;
   64538: out<=0;
   64539: out<=1;
   64540: out<=1;
   64541: out<=1;
   64542: out<=0;
   64543: out<=0;
   64544: out<=1;
   64545: out<=1;
   64546: out<=0;
   64547: out<=0;
   64548: out<=0;
   64549: out<=1;
   64550: out<=0;
   64551: out<=1;
   64552: out<=0;
   64553: out<=1;
   64554: out<=1;
   64555: out<=0;
   64556: out<=1;
   64557: out<=1;
   64558: out<=1;
   64559: out<=1;
   64560: out<=0;
   64561: out<=1;
   64562: out<=0;
   64563: out<=1;
   64564: out<=0;
   64565: out<=0;
   64566: out<=1;
   64567: out<=1;
   64568: out<=0;
   64569: out<=0;
   64570: out<=0;
   64571: out<=0;
   64572: out<=0;
   64573: out<=1;
   64574: out<=1;
   64575: out<=0;
   64576: out<=0;
   64577: out<=1;
   64578: out<=1;
   64579: out<=0;
   64580: out<=0;
   64581: out<=0;
   64582: out<=0;
   64583: out<=0;
   64584: out<=1;
   64585: out<=1;
   64586: out<=0;
   64587: out<=0;
   64588: out<=1;
   64589: out<=0;
   64590: out<=1;
   64591: out<=0;
   64592: out<=0;
   64593: out<=0;
   64594: out<=0;
   64595: out<=0;
   64596: out<=1;
   64597: out<=0;
   64598: out<=0;
   64599: out<=1;
   64600: out<=0;
   64601: out<=1;
   64602: out<=0;
   64603: out<=1;
   64604: out<=1;
   64605: out<=1;
   64606: out<=0;
   64607: out<=0;
   64608: out<=1;
   64609: out<=1;
   64610: out<=0;
   64611: out<=0;
   64612: out<=0;
   64613: out<=1;
   64614: out<=0;
   64615: out<=1;
   64616: out<=0;
   64617: out<=1;
   64618: out<=1;
   64619: out<=0;
   64620: out<=1;
   64621: out<=1;
   64622: out<=1;
   64623: out<=1;
   64624: out<=1;
   64625: out<=0;
   64626: out<=1;
   64627: out<=0;
   64628: out<=1;
   64629: out<=1;
   64630: out<=0;
   64631: out<=0;
   64632: out<=1;
   64633: out<=1;
   64634: out<=1;
   64635: out<=1;
   64636: out<=1;
   64637: out<=0;
   64638: out<=0;
   64639: out<=1;
   64640: out<=1;
   64641: out<=0;
   64642: out<=0;
   64643: out<=1;
   64644: out<=1;
   64645: out<=1;
   64646: out<=1;
   64647: out<=1;
   64648: out<=0;
   64649: out<=0;
   64650: out<=1;
   64651: out<=1;
   64652: out<=0;
   64653: out<=1;
   64654: out<=0;
   64655: out<=1;
   64656: out<=1;
   64657: out<=1;
   64658: out<=1;
   64659: out<=1;
   64660: out<=0;
   64661: out<=1;
   64662: out<=1;
   64663: out<=0;
   64664: out<=1;
   64665: out<=0;
   64666: out<=1;
   64667: out<=0;
   64668: out<=0;
   64669: out<=0;
   64670: out<=1;
   64671: out<=1;
   64672: out<=1;
   64673: out<=1;
   64674: out<=0;
   64675: out<=0;
   64676: out<=0;
   64677: out<=1;
   64678: out<=0;
   64679: out<=1;
   64680: out<=0;
   64681: out<=1;
   64682: out<=1;
   64683: out<=0;
   64684: out<=1;
   64685: out<=1;
   64686: out<=1;
   64687: out<=1;
   64688: out<=1;
   64689: out<=0;
   64690: out<=1;
   64691: out<=0;
   64692: out<=1;
   64693: out<=1;
   64694: out<=0;
   64695: out<=0;
   64696: out<=1;
   64697: out<=1;
   64698: out<=1;
   64699: out<=1;
   64700: out<=1;
   64701: out<=0;
   64702: out<=0;
   64703: out<=1;
   64704: out<=0;
   64705: out<=1;
   64706: out<=1;
   64707: out<=0;
   64708: out<=0;
   64709: out<=0;
   64710: out<=0;
   64711: out<=0;
   64712: out<=1;
   64713: out<=1;
   64714: out<=0;
   64715: out<=0;
   64716: out<=1;
   64717: out<=0;
   64718: out<=1;
   64719: out<=0;
   64720: out<=1;
   64721: out<=1;
   64722: out<=1;
   64723: out<=1;
   64724: out<=0;
   64725: out<=1;
   64726: out<=1;
   64727: out<=0;
   64728: out<=1;
   64729: out<=0;
   64730: out<=1;
   64731: out<=0;
   64732: out<=0;
   64733: out<=0;
   64734: out<=1;
   64735: out<=1;
   64736: out<=1;
   64737: out<=1;
   64738: out<=0;
   64739: out<=0;
   64740: out<=0;
   64741: out<=1;
   64742: out<=0;
   64743: out<=1;
   64744: out<=0;
   64745: out<=1;
   64746: out<=1;
   64747: out<=0;
   64748: out<=1;
   64749: out<=1;
   64750: out<=1;
   64751: out<=1;
   64752: out<=0;
   64753: out<=1;
   64754: out<=0;
   64755: out<=1;
   64756: out<=0;
   64757: out<=0;
   64758: out<=1;
   64759: out<=1;
   64760: out<=0;
   64761: out<=0;
   64762: out<=0;
   64763: out<=0;
   64764: out<=0;
   64765: out<=1;
   64766: out<=1;
   64767: out<=0;
   64768: out<=0;
   64769: out<=0;
   64770: out<=0;
   64771: out<=0;
   64772: out<=1;
   64773: out<=0;
   64774: out<=0;
   64775: out<=1;
   64776: out<=0;
   64777: out<=1;
   64778: out<=0;
   64779: out<=1;
   64780: out<=1;
   64781: out<=1;
   64782: out<=0;
   64783: out<=0;
   64784: out<=0;
   64785: out<=1;
   64786: out<=1;
   64787: out<=0;
   64788: out<=0;
   64789: out<=0;
   64790: out<=0;
   64791: out<=0;
   64792: out<=1;
   64793: out<=1;
   64794: out<=0;
   64795: out<=0;
   64796: out<=1;
   64797: out<=0;
   64798: out<=1;
   64799: out<=0;
   64800: out<=1;
   64801: out<=0;
   64802: out<=1;
   64803: out<=0;
   64804: out<=1;
   64805: out<=1;
   64806: out<=0;
   64807: out<=0;
   64808: out<=1;
   64809: out<=1;
   64810: out<=1;
   64811: out<=1;
   64812: out<=1;
   64813: out<=0;
   64814: out<=0;
   64815: out<=1;
   64816: out<=1;
   64817: out<=1;
   64818: out<=0;
   64819: out<=0;
   64820: out<=0;
   64821: out<=1;
   64822: out<=0;
   64823: out<=1;
   64824: out<=0;
   64825: out<=1;
   64826: out<=1;
   64827: out<=0;
   64828: out<=1;
   64829: out<=1;
   64830: out<=1;
   64831: out<=1;
   64832: out<=0;
   64833: out<=0;
   64834: out<=0;
   64835: out<=0;
   64836: out<=1;
   64837: out<=0;
   64838: out<=0;
   64839: out<=1;
   64840: out<=0;
   64841: out<=1;
   64842: out<=0;
   64843: out<=1;
   64844: out<=1;
   64845: out<=1;
   64846: out<=0;
   64847: out<=0;
   64848: out<=1;
   64849: out<=0;
   64850: out<=0;
   64851: out<=1;
   64852: out<=1;
   64853: out<=1;
   64854: out<=1;
   64855: out<=1;
   64856: out<=0;
   64857: out<=0;
   64858: out<=1;
   64859: out<=1;
   64860: out<=0;
   64861: out<=1;
   64862: out<=0;
   64863: out<=1;
   64864: out<=0;
   64865: out<=1;
   64866: out<=0;
   64867: out<=1;
   64868: out<=0;
   64869: out<=0;
   64870: out<=1;
   64871: out<=1;
   64872: out<=0;
   64873: out<=0;
   64874: out<=0;
   64875: out<=0;
   64876: out<=0;
   64877: out<=1;
   64878: out<=1;
   64879: out<=0;
   64880: out<=1;
   64881: out<=1;
   64882: out<=0;
   64883: out<=0;
   64884: out<=0;
   64885: out<=1;
   64886: out<=0;
   64887: out<=1;
   64888: out<=0;
   64889: out<=1;
   64890: out<=1;
   64891: out<=0;
   64892: out<=1;
   64893: out<=1;
   64894: out<=1;
   64895: out<=1;
   64896: out<=1;
   64897: out<=1;
   64898: out<=1;
   64899: out<=1;
   64900: out<=0;
   64901: out<=1;
   64902: out<=1;
   64903: out<=0;
   64904: out<=1;
   64905: out<=0;
   64906: out<=1;
   64907: out<=0;
   64908: out<=0;
   64909: out<=0;
   64910: out<=1;
   64911: out<=1;
   64912: out<=0;
   64913: out<=1;
   64914: out<=1;
   64915: out<=0;
   64916: out<=0;
   64917: out<=0;
   64918: out<=0;
   64919: out<=0;
   64920: out<=1;
   64921: out<=1;
   64922: out<=0;
   64923: out<=0;
   64924: out<=1;
   64925: out<=0;
   64926: out<=1;
   64927: out<=0;
   64928: out<=0;
   64929: out<=1;
   64930: out<=0;
   64931: out<=1;
   64932: out<=0;
   64933: out<=0;
   64934: out<=1;
   64935: out<=1;
   64936: out<=0;
   64937: out<=0;
   64938: out<=0;
   64939: out<=0;
   64940: out<=0;
   64941: out<=1;
   64942: out<=1;
   64943: out<=0;
   64944: out<=1;
   64945: out<=1;
   64946: out<=0;
   64947: out<=0;
   64948: out<=0;
   64949: out<=1;
   64950: out<=0;
   64951: out<=1;
   64952: out<=0;
   64953: out<=1;
   64954: out<=1;
   64955: out<=0;
   64956: out<=1;
   64957: out<=1;
   64958: out<=1;
   64959: out<=1;
   64960: out<=1;
   64961: out<=1;
   64962: out<=1;
   64963: out<=1;
   64964: out<=0;
   64965: out<=1;
   64966: out<=1;
   64967: out<=0;
   64968: out<=1;
   64969: out<=0;
   64970: out<=1;
   64971: out<=0;
   64972: out<=0;
   64973: out<=0;
   64974: out<=1;
   64975: out<=1;
   64976: out<=1;
   64977: out<=0;
   64978: out<=0;
   64979: out<=1;
   64980: out<=1;
   64981: out<=1;
   64982: out<=1;
   64983: out<=1;
   64984: out<=0;
   64985: out<=0;
   64986: out<=1;
   64987: out<=1;
   64988: out<=0;
   64989: out<=1;
   64990: out<=0;
   64991: out<=1;
   64992: out<=1;
   64993: out<=0;
   64994: out<=1;
   64995: out<=0;
   64996: out<=1;
   64997: out<=1;
   64998: out<=0;
   64999: out<=0;
   65000: out<=1;
   65001: out<=1;
   65002: out<=1;
   65003: out<=1;
   65004: out<=1;
   65005: out<=0;
   65006: out<=0;
   65007: out<=1;
   65008: out<=1;
   65009: out<=1;
   65010: out<=0;
   65011: out<=0;
   65012: out<=0;
   65013: out<=1;
   65014: out<=0;
   65015: out<=1;
   65016: out<=0;
   65017: out<=1;
   65018: out<=1;
   65019: out<=0;
   65020: out<=1;
   65021: out<=1;
   65022: out<=1;
   65023: out<=1;
   65024: out<=1;
   65025: out<=1;
   65026: out<=0;
   65027: out<=0;
   65028: out<=0;
   65029: out<=1;
   65030: out<=0;
   65031: out<=1;
   65032: out<=0;
   65033: out<=1;
   65034: out<=1;
   65035: out<=0;
   65036: out<=1;
   65037: out<=1;
   65038: out<=1;
   65039: out<=1;
   65040: out<=1;
   65041: out<=0;
   65042: out<=1;
   65043: out<=0;
   65044: out<=1;
   65045: out<=1;
   65046: out<=0;
   65047: out<=0;
   65048: out<=1;
   65049: out<=1;
   65050: out<=1;
   65051: out<=1;
   65052: out<=1;
   65053: out<=0;
   65054: out<=0;
   65055: out<=1;
   65056: out<=1;
   65057: out<=0;
   65058: out<=0;
   65059: out<=1;
   65060: out<=1;
   65061: out<=1;
   65062: out<=1;
   65063: out<=1;
   65064: out<=0;
   65065: out<=0;
   65066: out<=1;
   65067: out<=1;
   65068: out<=0;
   65069: out<=1;
   65070: out<=0;
   65071: out<=1;
   65072: out<=1;
   65073: out<=1;
   65074: out<=1;
   65075: out<=1;
   65076: out<=0;
   65077: out<=1;
   65078: out<=1;
   65079: out<=0;
   65080: out<=1;
   65081: out<=0;
   65082: out<=1;
   65083: out<=0;
   65084: out<=0;
   65085: out<=0;
   65086: out<=1;
   65087: out<=1;
   65088: out<=1;
   65089: out<=1;
   65090: out<=0;
   65091: out<=0;
   65092: out<=0;
   65093: out<=1;
   65094: out<=0;
   65095: out<=1;
   65096: out<=0;
   65097: out<=1;
   65098: out<=1;
   65099: out<=0;
   65100: out<=1;
   65101: out<=1;
   65102: out<=1;
   65103: out<=1;
   65104: out<=0;
   65105: out<=1;
   65106: out<=0;
   65107: out<=1;
   65108: out<=0;
   65109: out<=0;
   65110: out<=1;
   65111: out<=1;
   65112: out<=0;
   65113: out<=0;
   65114: out<=0;
   65115: out<=0;
   65116: out<=0;
   65117: out<=1;
   65118: out<=1;
   65119: out<=0;
   65120: out<=0;
   65121: out<=1;
   65122: out<=1;
   65123: out<=0;
   65124: out<=0;
   65125: out<=0;
   65126: out<=0;
   65127: out<=0;
   65128: out<=1;
   65129: out<=1;
   65130: out<=0;
   65131: out<=0;
   65132: out<=1;
   65133: out<=0;
   65134: out<=1;
   65135: out<=0;
   65136: out<=1;
   65137: out<=1;
   65138: out<=1;
   65139: out<=1;
   65140: out<=0;
   65141: out<=1;
   65142: out<=1;
   65143: out<=0;
   65144: out<=1;
   65145: out<=0;
   65146: out<=1;
   65147: out<=0;
   65148: out<=0;
   65149: out<=0;
   65150: out<=1;
   65151: out<=1;
   65152: out<=1;
   65153: out<=1;
   65154: out<=0;
   65155: out<=0;
   65156: out<=0;
   65157: out<=1;
   65158: out<=0;
   65159: out<=1;
   65160: out<=0;
   65161: out<=1;
   65162: out<=1;
   65163: out<=0;
   65164: out<=1;
   65165: out<=1;
   65166: out<=1;
   65167: out<=1;
   65168: out<=0;
   65169: out<=1;
   65170: out<=0;
   65171: out<=1;
   65172: out<=0;
   65173: out<=0;
   65174: out<=1;
   65175: out<=1;
   65176: out<=0;
   65177: out<=0;
   65178: out<=0;
   65179: out<=0;
   65180: out<=0;
   65181: out<=1;
   65182: out<=1;
   65183: out<=0;
   65184: out<=1;
   65185: out<=0;
   65186: out<=0;
   65187: out<=1;
   65188: out<=1;
   65189: out<=1;
   65190: out<=1;
   65191: out<=1;
   65192: out<=0;
   65193: out<=0;
   65194: out<=1;
   65195: out<=1;
   65196: out<=0;
   65197: out<=1;
   65198: out<=0;
   65199: out<=1;
   65200: out<=0;
   65201: out<=0;
   65202: out<=0;
   65203: out<=0;
   65204: out<=1;
   65205: out<=0;
   65206: out<=0;
   65207: out<=1;
   65208: out<=0;
   65209: out<=1;
   65210: out<=0;
   65211: out<=1;
   65212: out<=1;
   65213: out<=1;
   65214: out<=0;
   65215: out<=0;
   65216: out<=1;
   65217: out<=1;
   65218: out<=0;
   65219: out<=0;
   65220: out<=0;
   65221: out<=1;
   65222: out<=0;
   65223: out<=1;
   65224: out<=0;
   65225: out<=1;
   65226: out<=1;
   65227: out<=0;
   65228: out<=1;
   65229: out<=1;
   65230: out<=1;
   65231: out<=1;
   65232: out<=1;
   65233: out<=0;
   65234: out<=1;
   65235: out<=0;
   65236: out<=1;
   65237: out<=1;
   65238: out<=0;
   65239: out<=0;
   65240: out<=1;
   65241: out<=1;
   65242: out<=1;
   65243: out<=1;
   65244: out<=1;
   65245: out<=0;
   65246: out<=0;
   65247: out<=1;
   65248: out<=0;
   65249: out<=1;
   65250: out<=1;
   65251: out<=0;
   65252: out<=0;
   65253: out<=0;
   65254: out<=0;
   65255: out<=0;
   65256: out<=1;
   65257: out<=1;
   65258: out<=0;
   65259: out<=0;
   65260: out<=1;
   65261: out<=0;
   65262: out<=1;
   65263: out<=0;
   65264: out<=0;
   65265: out<=0;
   65266: out<=0;
   65267: out<=0;
   65268: out<=1;
   65269: out<=0;
   65270: out<=0;
   65271: out<=1;
   65272: out<=0;
   65273: out<=1;
   65274: out<=0;
   65275: out<=1;
   65276: out<=1;
   65277: out<=1;
   65278: out<=0;
   65279: out<=0;
   65280: out<=0;
   65281: out<=1;
   65282: out<=0;
   65283: out<=1;
   65284: out<=0;
   65285: out<=0;
   65286: out<=1;
   65287: out<=1;
   65288: out<=0;
   65289: out<=0;
   65290: out<=0;
   65291: out<=0;
   65292: out<=0;
   65293: out<=1;
   65294: out<=1;
   65295: out<=0;
   65296: out<=1;
   65297: out<=1;
   65298: out<=0;
   65299: out<=0;
   65300: out<=0;
   65301: out<=1;
   65302: out<=0;
   65303: out<=1;
   65304: out<=0;
   65305: out<=1;
   65306: out<=1;
   65307: out<=0;
   65308: out<=1;
   65309: out<=1;
   65310: out<=1;
   65311: out<=1;
   65312: out<=1;
   65313: out<=1;
   65314: out<=1;
   65315: out<=1;
   65316: out<=0;
   65317: out<=1;
   65318: out<=1;
   65319: out<=0;
   65320: out<=1;
   65321: out<=0;
   65322: out<=1;
   65323: out<=0;
   65324: out<=0;
   65325: out<=0;
   65326: out<=1;
   65327: out<=1;
   65328: out<=0;
   65329: out<=1;
   65330: out<=1;
   65331: out<=0;
   65332: out<=0;
   65333: out<=0;
   65334: out<=0;
   65335: out<=0;
   65336: out<=1;
   65337: out<=1;
   65338: out<=0;
   65339: out<=0;
   65340: out<=1;
   65341: out<=0;
   65342: out<=1;
   65343: out<=0;
   65344: out<=1;
   65345: out<=0;
   65346: out<=1;
   65347: out<=0;
   65348: out<=1;
   65349: out<=1;
   65350: out<=0;
   65351: out<=0;
   65352: out<=1;
   65353: out<=1;
   65354: out<=1;
   65355: out<=1;
   65356: out<=1;
   65357: out<=0;
   65358: out<=0;
   65359: out<=1;
   65360: out<=1;
   65361: out<=1;
   65362: out<=0;
   65363: out<=0;
   65364: out<=0;
   65365: out<=1;
   65366: out<=0;
   65367: out<=1;
   65368: out<=0;
   65369: out<=1;
   65370: out<=1;
   65371: out<=0;
   65372: out<=1;
   65373: out<=1;
   65374: out<=1;
   65375: out<=1;
   65376: out<=1;
   65377: out<=1;
   65378: out<=1;
   65379: out<=1;
   65380: out<=0;
   65381: out<=1;
   65382: out<=1;
   65383: out<=0;
   65384: out<=1;
   65385: out<=0;
   65386: out<=1;
   65387: out<=0;
   65388: out<=0;
   65389: out<=0;
   65390: out<=1;
   65391: out<=1;
   65392: out<=1;
   65393: out<=0;
   65394: out<=0;
   65395: out<=1;
   65396: out<=1;
   65397: out<=1;
   65398: out<=1;
   65399: out<=1;
   65400: out<=0;
   65401: out<=0;
   65402: out<=1;
   65403: out<=1;
   65404: out<=0;
   65405: out<=1;
   65406: out<=0;
   65407: out<=1;
   65408: out<=1;
   65409: out<=0;
   65410: out<=1;
   65411: out<=0;
   65412: out<=1;
   65413: out<=1;
   65414: out<=0;
   65415: out<=0;
   65416: out<=1;
   65417: out<=1;
   65418: out<=1;
   65419: out<=1;
   65420: out<=1;
   65421: out<=0;
   65422: out<=0;
   65423: out<=1;
   65424: out<=1;
   65425: out<=1;
   65426: out<=0;
   65427: out<=0;
   65428: out<=0;
   65429: out<=1;
   65430: out<=0;
   65431: out<=1;
   65432: out<=0;
   65433: out<=1;
   65434: out<=1;
   65435: out<=0;
   65436: out<=1;
   65437: out<=1;
   65438: out<=1;
   65439: out<=1;
   65440: out<=0;
   65441: out<=0;
   65442: out<=0;
   65443: out<=0;
   65444: out<=1;
   65445: out<=0;
   65446: out<=0;
   65447: out<=1;
   65448: out<=0;
   65449: out<=1;
   65450: out<=0;
   65451: out<=1;
   65452: out<=1;
   65453: out<=1;
   65454: out<=0;
   65455: out<=0;
   65456: out<=0;
   65457: out<=1;
   65458: out<=1;
   65459: out<=0;
   65460: out<=0;
   65461: out<=0;
   65462: out<=0;
   65463: out<=0;
   65464: out<=1;
   65465: out<=1;
   65466: out<=0;
   65467: out<=0;
   65468: out<=1;
   65469: out<=0;
   65470: out<=1;
   65471: out<=0;
   65472: out<=0;
   65473: out<=1;
   65474: out<=0;
   65475: out<=1;
   65476: out<=0;
   65477: out<=0;
   65478: out<=1;
   65479: out<=1;
   65480: out<=0;
   65481: out<=0;
   65482: out<=0;
   65483: out<=0;
   65484: out<=0;
   65485: out<=1;
   65486: out<=1;
   65487: out<=0;
   65488: out<=1;
   65489: out<=1;
   65490: out<=0;
   65491: out<=0;
   65492: out<=0;
   65493: out<=1;
   65494: out<=0;
   65495: out<=1;
   65496: out<=0;
   65497: out<=1;
   65498: out<=1;
   65499: out<=0;
   65500: out<=1;
   65501: out<=1;
   65502: out<=1;
   65503: out<=1;
   65504: out<=0;
   65505: out<=0;
   65506: out<=0;
   65507: out<=0;
   65508: out<=1;
   65509: out<=0;
   65510: out<=0;
   65511: out<=1;
   65512: out<=0;
   65513: out<=1;
   65514: out<=0;
   65515: out<=1;
   65516: out<=1;
   65517: out<=1;
   65518: out<=0;
   65519: out<=0;
   65520: out<=1;
   65521: out<=0;
   65522: out<=0;
   65523: out<=1;
   65524: out<=1;
   65525: out<=1;
   65526: out<=1;
   65527: out<=1;
   65528: out<=0;
   65529: out<=0;
   65530: out<=1;
   65531: out<=1;
   65532: out<=0;
   65533: out<=1;
   65534: out<=0;
   65535: out<=1;
 endcase
end
endmodule
