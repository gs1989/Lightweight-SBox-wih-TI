module STI4_R2_191(in,out);
  input[7:0] in;
  output out;
  reg out;
  always@(in)
  begin
    case(in)
   0: out<=0;
   1: out<=0;
   2: out<=1;
   3: out<=0;
   4: out<=1;
   5: out<=0;
   6: out<=0;
   7: out<=0;
   8: out<=1;
   9: out<=1;
   10: out<=1;
   11: out<=0;
   12: out<=1;
   13: out<=0;
   14: out<=1;
   15: out<=1;
   16: out<=0;
   17: out<=0;
   18: out<=0;
   19: out<=1;
   20: out<=0;
   21: out<=1;
   22: out<=0;
   23: out<=0;
   24: out<=1;
   25: out<=1;
   26: out<=0;
   27: out<=1;
   28: out<=0;
   29: out<=1;
   30: out<=1;
   31: out<=1;
   32: out<=0;
   33: out<=1;
   34: out<=1;
   35: out<=1;
   36: out<=1;
   37: out<=1;
   38: out<=0;
   39: out<=1;
   40: out<=0;
   41: out<=1;
   42: out<=0;
   43: out<=0;
   44: out<=0;
   45: out<=0;
   46: out<=0;
   47: out<=1;
   48: out<=0;
   49: out<=1;
   50: out<=0;
   51: out<=0;
   52: out<=0;
   53: out<=0;
   54: out<=0;
   55: out<=1;
   56: out<=0;
   57: out<=1;
   58: out<=1;
   59: out<=1;
   60: out<=1;
   61: out<=1;
   62: out<=0;
   63: out<=1;
   64: out<=0;
   65: out<=1;
   66: out<=1;
   67: out<=1;
   68: out<=1;
   69: out<=1;
   70: out<=0;
   71: out<=1;
   72: out<=0;
   73: out<=1;
   74: out<=0;
   75: out<=0;
   76: out<=0;
   77: out<=0;
   78: out<=0;
   79: out<=1;
   80: out<=0;
   81: out<=1;
   82: out<=0;
   83: out<=0;
   84: out<=0;
   85: out<=0;
   86: out<=0;
   87: out<=1;
   88: out<=0;
   89: out<=1;
   90: out<=1;
   91: out<=1;
   92: out<=1;
   93: out<=1;
   94: out<=0;
   95: out<=1;
   96: out<=0;
   97: out<=0;
   98: out<=1;
   99: out<=0;
   100: out<=1;
   101: out<=0;
   102: out<=0;
   103: out<=0;
   104: out<=1;
   105: out<=1;
   106: out<=1;
   107: out<=0;
   108: out<=1;
   109: out<=0;
   110: out<=1;
   111: out<=1;
   112: out<=0;
   113: out<=0;
   114: out<=0;
   115: out<=1;
   116: out<=0;
   117: out<=1;
   118: out<=0;
   119: out<=0;
   120: out<=1;
   121: out<=1;
   122: out<=0;
   123: out<=1;
   124: out<=0;
   125: out<=1;
   126: out<=1;
   127: out<=1;
   128: out<=0;
   129: out<=0;
   130: out<=0;
   131: out<=1;
   132: out<=0;
   133: out<=1;
   134: out<=0;
   135: out<=0;
   136: out<=1;
   137: out<=1;
   138: out<=0;
   139: out<=1;
   140: out<=0;
   141: out<=1;
   142: out<=1;
   143: out<=1;
   144: out<=0;
   145: out<=0;
   146: out<=1;
   147: out<=0;
   148: out<=1;
   149: out<=0;
   150: out<=0;
   151: out<=0;
   152: out<=1;
   153: out<=1;
   154: out<=1;
   155: out<=0;
   156: out<=1;
   157: out<=0;
   158: out<=1;
   159: out<=1;
   160: out<=0;
   161: out<=1;
   162: out<=0;
   163: out<=0;
   164: out<=0;
   165: out<=0;
   166: out<=0;
   167: out<=1;
   168: out<=0;
   169: out<=1;
   170: out<=1;
   171: out<=1;
   172: out<=1;
   173: out<=1;
   174: out<=0;
   175: out<=1;
   176: out<=0;
   177: out<=1;
   178: out<=1;
   179: out<=1;
   180: out<=1;
   181: out<=1;
   182: out<=0;
   183: out<=1;
   184: out<=0;
   185: out<=1;
   186: out<=0;
   187: out<=0;
   188: out<=0;
   189: out<=0;
   190: out<=0;
   191: out<=1;
   192: out<=0;
   193: out<=1;
   194: out<=0;
   195: out<=0;
   196: out<=0;
   197: out<=0;
   198: out<=0;
   199: out<=1;
   200: out<=0;
   201: out<=1;
   202: out<=1;
   203: out<=1;
   204: out<=1;
   205: out<=1;
   206: out<=0;
   207: out<=1;
   208: out<=0;
   209: out<=1;
   210: out<=1;
   211: out<=1;
   212: out<=1;
   213: out<=1;
   214: out<=0;
   215: out<=1;
   216: out<=0;
   217: out<=1;
   218: out<=0;
   219: out<=0;
   220: out<=0;
   221: out<=0;
   222: out<=0;
   223: out<=1;
   224: out<=0;
   225: out<=0;
   226: out<=0;
   227: out<=1;
   228: out<=0;
   229: out<=1;
   230: out<=0;
   231: out<=0;
   232: out<=1;
   233: out<=1;
   234: out<=0;
   235: out<=1;
   236: out<=0;
   237: out<=1;
   238: out<=1;
   239: out<=1;
   240: out<=0;
   241: out<=0;
   242: out<=1;
   243: out<=0;
   244: out<=1;
   245: out<=0;
   246: out<=0;
   247: out<=0;
   248: out<=1;
   249: out<=1;
   250: out<=1;
   251: out<=0;
   252: out<=1;
   253: out<=0;
   254: out<=1;
   255: out<=1;
 endcase
end
endmodule
